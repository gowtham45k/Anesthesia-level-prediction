��
      �yellowbrick.regressor.residuals��ResidualsPlot���)��}�(�force_model���	estimator��sklearn.linear_model._base��LinearRegression���)��}�(�fit_intercept���copy_X���n_jobs�N�positive���n_features_in_�K	�coef_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK	��h�dtype����f8�����R�(K�<�NNNJ����J����K t�b�CHF�j��)Q?ۛ�j��j?^�]��?>�'R?]�9�h?�Dm�0����I��W?��a
�i�B�&:픎?�t�b�rank_�K	�	singular_�hhK ��h��R�(KK	��h!�CH��0�y�@��#�>Zv@ɛ�M^Ri@����3b@MI;��/T@خ:�N@3�I��{C@�W��i'@�a��w�&@�t�b�
intercept_�h�scalar���h!CvӕW��?���R��_sklearn_version��1.4.1.post1�ub�	is_fitted��auto��name�h�_wrapped�h
�_ax��matplotlib.axes._axes��Axes���)��}�(�_stale���stale_callback�N�_axes�h>�figure��matplotlib.figure��Figure���)��}�(h@�hANhChG�
_transform�N�_transformSet���_visible���	_animated���_alpha�N�clipbox�N�	_clippath�N�_clipon���_label�� ��_picker�N�_rasterized���_agg_filter�N�
_mouseover���
_callbacks��matplotlib.cbook��CallbackRegistry���)��}�(�_signals�]��pchanged�a�exception_handler�hX�_exception_printer����	callbacks�}��_cid_gen�K �_func_cid_map�N�_pickled_cids���ub�_remove_method�N�_url�N�_gid�N�_snap�N�_sketch�N�_path_effects�]��_sticky_edges��matplotlib.artist��_XYPair���]�]������
_in_layout���	_suptitle�N�
_supxlabel�N�
_supylabel�N�_align_label_groups�}�(�x�hX�Grouper���)��}��_mapping�}�sb�y�h�)��}�h�}�sbu�
_localaxes�]�(h>h=)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhi�builtins��getattr���hG�delaxes���R�hjNhkNhlNhmNhnhohphs]�]�����hx��	_position��matplotlib.transforms��Bbox���)��}�(�_parents�}�����Hh��TransformedBbox���)��}�(h�}��P��Hh��BboxTransformTo���)��}�(h�}�(����Hh��CompositeGenericTransform���)��}�(�
input_dims�K�output_dims�Kh�}��О�Hh�)��}�(h�Kh�Kh�}�(����Hh��BlendedGenericTransform���)��}�(h�}�(���Hh�)��}�(h�Kh�Kh�}��_invalid�K�_shorthand_name�hR�_a�h��_b�h��ScaledTranslation���)��}�(h�}����Hh�sh�K h�hR�	_inverted�N�_t�K G���8�9���_scale_trans�h��Affine2D���)��}�(h�}�(�����Hh�)��}�(h�}��P���Hh�)��}�(h�}�(��-��Hh�)��}�(h�}���
�Hh�)��}�(h�}�(��+��Hh�)��}�(h�Kh�Kh�}���[�Hh�)��}�(h�Kh�Kh�}�(�PzS�Hh�)��}�(h�}�(�PV�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��PV�Hh�sh�K h�hRh�Nh�K G���8�9��h�hό_mtx�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bubub�Pn��Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��Pn��Hh�sh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nubub���Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}����Hh�sh�K h�hRh�Nh�K G���8�9��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bubub�p�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��p�Hj	  sh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nubub�H�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��H�Hj  sh�Kh�hRh�Nh�K G��-��-�؆�h�h�h�Nubub�Ќ�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}��Ќ�Hj  sh�Kh�hRh�Nh�K G?�-��-�؆�h�h�h�Nubub��^�Hh��TransformedPath���)��}�(h�}�h�Kh�hR�_path��matplotlib.path��Path���)��}�(�	_vertices�hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�b�_codes�N�_interpolation_steps�K��_simplify_threshold�G?�q�q�֌_should_simplify���	_readonly��ubhIh�_transformed_path�j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ub�_transformed_points�j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��!�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�3!�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P� �Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P""�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?      �?              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P)"�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        @       @              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P`�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       @      @              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P� �Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       @      @              �?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIh�j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ububuh�Kh�hR�_x�h�_y�hی_affine�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CHŠk�.p@        
�J�\�             xz@9��8��I@                      �?�t�bubub��
�Hh�)��}�(h�}�(��Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}���Hj�  sh�K h�hRh�Nh�G���8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#�              �?                              �?�t�bubub�	�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}��	�Hj�  sh�Kh�hRh�Nh�G?��8�9K ��h�h�h�Nubub��#�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}���#�Hj�  sh�K h�hRh�Nh�G���8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#�              �?                              �?�t�bubub�'�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}��'�Hj�  sh�Kh�hRh�Nh�G?��8�9K ��h�h�h�Nubub�P��Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}��P��Hj�  sh�Kh�hRh�Nh�G��-��-��K ��h�h�h�Nubub�п�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j�  h�h�)��}�(h�}��п�Hj�  sh�Kh�hRh�Nh�G?�-��-��K ��h�h�h�Nubub�����Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubub����Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�433333㿔t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��3�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ٿ������ٿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub����Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ɿ������ɿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��8�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j,  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P��Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  j;  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j;  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�Pn��Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  jJ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jJ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P� �Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�?433333�?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj�  j5  j&  )��}�(j)  jY  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jY  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ububuh�Kh�hRj�  h�j�  h�j�  h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@        ���@;t@����l�o@                      �?�t�bububuh�Kh�hRh�h��TransformWrapper���)��}�(h�}�(�P[c�Hh�)��}�(h�}��P�
�Hh��BboxTransformFrom���)��}�(h�}���+��Hh�sh�K h�hRh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH��l%��?        �Ԓ.�p�?        �v����?����p�                      �?�t�bub�_boxin�jo  h�hhK ��h��R�(KKK��h!�CH�!��>�?        ��d*R�ֿ        ��tSau�?�S�Ġ��?                      �?�t�bubsh�K h�hR�_bbox�h�)��}�(h�}��P[c�Hjo  sh�K h�hR�_points�hhK ��h��R�(KKK��h!�C �Ԓ.�p�?����p俲[8^@�J�Qv��?�t�b�_minpos�hhK ��h��R�(KK��h!�C      �      ��t�b�_ignore���_points_orig�hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjl  j�  hhK ��h��R�(KKK��h!�C �Ԓ.�p�?����p俲[8^@�J�Qv��?�t�bub��[�Hh�uh�K h�hR�_child�h��BlendedAffine2D���)��}�(h�}����Hjl  sh�K h�hRj�  h��IdentityTransform���)��}�(h�}��P��Hj�  sh�Kh�hRh�Nubj�  j�  )��}�(h�}��P��Hj�  sh�Kh�hRh�Nubh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bub�	transform�h�j�  j�  ��R��transform_affine�h�j�  j�  ��R��transform_non_affine�h�j�  j�  ��R��transform_path�h�j�  j�  ��R��transform_path_affine�h�j�  j�  ��R��transform_path_non_affine�h�j�  j�  ��R��
get_affine�h�j�  j�  ��R��inverted�h�j�  j�  ��R��
get_matrix�h�j�  j�  ��R�ubh�h�ubsh�Kh�hRh�jt  h�h�ub�PzS�Hh��
�Hj�  ��[S�Hj�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}���[S�Hj�  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@              �?                              �?�t�bub���i�Hj�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}����i�Hj�  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH     �@              Y@              �?                              �?�t�bub�Е��Hj�  )��}�(h�}�h�Kh�hRj�  j�  )��}�(h�}��Е��Hj�  sh�Kh�hRh�Nubj�  h�h�Nh�hhK ��h��R�(KKK��h!�CH      �?                             xz@9��8��I@                      �?�t�bub�PP��Hj�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}��PP��Hj  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@              �?                              �?�t�bub��1�Hh�)��}�(h�Kh�Kh�}��2�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��2�Hj  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���1�Hj  sh�Kh�hRh�h�)��}�(h�}��P1�Hj*  sh�Kh�hRh�N�_boxout�h�)��}�(h�}��0�Hj-  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P1�Hj*  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}�����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����HjR  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjO  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��HjO  sh�Kh�hRh�h�)��}�(h�}��Џ�Hjj  sh�Kh�hRh�Nj0  h�)��}�(h�}����Hjm  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��Џ�Hjj  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�  sh�Kh�hRh�h�)��}�(h�}�����Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�:�Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��:�Hj�  sh�Kh�hRh�h�)��}�(h�}��P7�Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}���:�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P7�Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}�����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��Hj  sh�Kh�hRh�h�)��}�(h�}����Hj9  sh�K h�hRh�Nj0  h�)��}�(h�}��P��Hj<  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj9  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}�����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����Hjf  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjc  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��Hjc  sh�Kh�hRh�h�)��}�(h�}��Й�Hj~  sh�Kh�hRh�Nj0  h�)��}�(h�}�����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��Й�Hj~  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�  sh�Kh�hRh�h�)��}�(h�}�����Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}�����Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�  sh�Kh�hRh�h�)��}�(h�}�����Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}�����Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Ђ�Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj#  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj   j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Ђ�Hj   sh�Kh�hRh�h�)��}�(h�}�����Hj;  sh�Kh�hRh�Nj0  h�)��}�(h�}����Hj>  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}�����Hj;  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����Hh�)��}�(h�Kh�Kh�}��І�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��І�Hjb  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj_  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����Hj_  sh�Kh�hRh�h�)��}�(h�}����Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��Є�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}�����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����Hj�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��Hj�  sh�Kh�hRh�h�)��}�(h�}��Љ�Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}�����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��Љ�Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�  sh�Kh�hRh�h�)��}�(h�}�����Hj
  sh�K h�hRh�Nj0  h�)��}�(h�}��P��Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����Hj
  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Б�Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj7  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj4  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Б�Hj4  sh�Kh�hRh�h�)��}�(h�}��P��HjO  sh�Kh�hRh�Nj0  h�)��}�(h�}����HjR  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P��HjO  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����Hh�)��}�(h�Kh�Kh�}��Е�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Е�Hjv  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjs  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����Hjs  sh�Kh�hRh�h�)��}�(h�}����Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}��Г�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}����Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�V�Hh�)��}�(h�Kh�Kh�}��b�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��b�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��V�Hj�  sh�Kh�hRh�h�)��}�(h�}���Q�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���l�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���Q�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�Hj�  sh�Kh�hRh�h�)��}�(h�}��P�Hj  sh�K h�hRh�Nj0  h�)��}�(h�}��P�Hj!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�h�)��}�(h�}�(����HjH  �P�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�jK  ub��+�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�jK  ubuh�K h�hRh�Nh�G        G?�UUUUUU��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?������ @                      �?�t�bubub�P�HjN  ��+�HjQ  ��Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj^  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj[  j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���Hj[  sh�Kh�hRh�h�)��}�(h�}���<�Hj|  sh�K h�hRh�Nj0  h�)��}�(h�}���%�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���<�Hj|  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ubuh�Kh�hRh�Nj0  h�h�hhK ��h��R�(KKK��h!�CH    �@        �qǱP@             xz@9��8��I@                      �?�t�bubsh�Kh�hRj�  h�)��}�(h�}���-��Hh�sh�K h�hRj�  hhK ��h��R�(KKK��h!�C       �?(\���(�?ffffff�?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIh�j�  hhK ��h��R�(KKK��h!�C �qǱP@9��8��I@�8��8�@�q�q�}@�t�bub����Hh�uh�Kh�hRh�Nj0  h�h�hhK ��h��R�(KKK��h!�CH      �@        �q�q�@�             0�@�q�q"�                      �?�t�bubsh�K h�hRj�  h�)��}�(h�}������Hh�sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                        @      @�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                        @      @�t�bubhIh�j�  hhK ��h��R�(KKK��h!�C                       �@     0�@�t�bub���	�Hh�P���Hh����Hh���R�Hj  ����Hj�  ��
�Hj�  ��$��Hj�  ���Hj�  �"�Hj  ���Hj  �Pah�Hj�  ����Hj�  �P���HhƊ��Hh�)��}�(h�}����Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nub�Po�Hh�)��}�(h�}����Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�K h�hRh�Nh�K G���8�9��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bub��q�Hh�)��}�(h�}�����Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G?��8�9��h�h�h�Nub����Hh�)��}�(h�}����Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�)��}�(h�}�(���Hj  �P��Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}��P��Hj  sh�K h�hRh�Nh�G?��8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#@              �?                              �?�t�bubub��I�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}���I�Hj  sh�Kh�hRh�Nh�G���8�9K ��h�h�h�Nubub��K�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}���K�Hj   sh�K h�hRh�Nh�G?��8�9K ��h�h�h�hhK ��h��R�(KKK��h!�CH      �?        �q�q#@              �?                              �?�t�bubub��"�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}���"�Hj-  sh�Kh�hRh�Nh�G��-��-��K ��h�h�h�Nubub�P&�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�j	  h�h�)��}�(h�}��P&�Hj4  sh�Kh�hRh�Nh�G?�-��-��K ��h�h�h�Nubub�P�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubj8  j&  )��}�(j)  jB  j0  Nj4  �j3  �j2  G?�q�q��j1  Kubub��!&�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�433333㿔t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jQ  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��&�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ٿ������ٿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j`  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�P��Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?������ɿ������ɿ�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  jo  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�Q'�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?                �t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j~  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�W'�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub�Px'�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?�������?�������?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubub��&�Hj  )��}�(h�}�h�Kh�hRj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?433333�?433333�?�t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubhIj	  j5  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ubj8  j&  )��}�(j)  j�  j0  Nj4  �j3  �j2  G?�q�q��j1  K�ububuh�Kh�hRj�  h�j�  h�j�  h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �8��8V�@        ���@;t@����l�o@                      �?�t�bububh�j  ubsh�Kh�hRh�Nh�G���8�9K ��h�h�h�Nub�P#�Hj  ���Hj  ����Hj#  �G4�Hh�)��}�(h�}�(���Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ub���Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ub�P��Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubuh�K h�hRh�Nh�G        G?�UUUUUU��h�h�h�hhK ��h��R�(KKK��h!�CH      �?                              �?������ @                      �?�t�bub����Hh�)��}�(h�}��m�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G��-��-�؆�h�h�h�Nub��o�Hh�)��}�(h�}��n�Hh�)��}�(h�Kh�Kh�}�h�Kh�hRh�h�h�j�  ubsh�Kh�hRh�Nh�K G?�-��-�؆�h�h�h�Nub�P$�Hj0  ��%�Hj7  �PT�HjK  uh�K h�hRh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH{�G�z�?                        {�G�z�?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      Y@                              Y@                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?�q�q#�                      �?�t�bubub���Hj�  ���Hj�  ����Hj�  �m�Hj�  �n�Hj�  uh�Kh�hRj�  h�j�  h�j�  h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CHn�d���@        �8��8V�@             xz@9��8��I@                      �?�t�bubub�P��Hj	  uh�Kh�hRh�jk  )��}�(h�}�(�Н�Hh�)��}�(h�}�����Hjs  )��}�(h�}�����Hh�sh�K h�hRh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH33333�F@                        �v����?����p�                      �?�t�bubj�  j�  h�hhK ��h��R�(KKK��h!�CH�����?               �        ��tSau�?�S�Ġ��?                      �?�t�bubsh�K h�hRj�  h�)��}�(h�}��Н�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C         ����p�33333�F@�J�Qv��?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C         ����p�33333�F@�J�Qv��?�t�bub�О�Hh�uh�K h�hRj�  j�  )��}�(h�}��С�Hj�  sh�K h�hRj�  j�  )��}�(h�}��R�Hj/	  sh�Kh�hRh�Nubj�  j�  )��}�(h�}��R�Hj/	  sh�Kh�hRh�Nubh�h�)��}�(h�}�h�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�j�  ubj�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�j�  h�j/	  j�  ��R�ubh�h�ubsh�Kh�hRh�j	  h�h�ub����Hh��P��Hj	  ��9l�Hj�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}���9l�HjS	  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �8��8V�@              �?                              �?�t�bub��Hj�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}���Hj_	  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �����_�@              �?                              �?�t�bub����Hj�  )��}�(h�}�h�Kh�hRj�  j�  )��}�(h�}�����Hjk	  sh�Kh�hRh�Nubj�  h�h�Nh�hhK ��h��R�(KKK��h!�CH      �?                             xz@�����?N@                      �?�t�bub�P��Hj�  )��}�(h�}�h�Kh�hRj�  h�j�  j�  )��}�(h�}��P��Hjw	  sh�Kh�hRh�Nubh�Nh�hhK ��h��R�(KKK��h!�CH      Y@        �����_�@              �?                              �?�t�bub���Hj�  ���Hj�  �P��Hj�  ��}�Hh�)��}�(h�Kh�Kh�}��P~�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P~�Hj�	  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�	  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���}�Hj�	  sh�Kh�hRh�h�)��}�(h�}���j�Hj�	  sh�Kh�hRh�Nj0  h�)��}�(h�}�����Hj�	  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���j�Hj�	  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��p�Hh�)��}�(h�Kh�Kh�}��q�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��q�Hj�	  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�	  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���p�Hj�	  sh�Kh�hRh�h�)��}�(h�}���j�Hj�	  sh�Kh�hRh�Nj0  h�)��}�(h�}���n�Hj�	  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���j�Hj�	  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pt�Hh�)��}�(h�Kh�Kh�}���t�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���t�Hj
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pt�Hj
  sh�Kh�hRh�h�)��}�(h�}���s�Hj
  sh�Kh�hRh�Nj0  h�)��}�(h�}���r�Hj
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���s�Hj
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�x�Hh�)��}�(h�Kh�Kh�}��Px�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Px�HjC
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj@
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��x�Hj@
  sh�Kh�hRh�h�)��}�(h�}���w�Hj[
  sh�Kh�hRh�Nj0  h�)��}�(h�}��Pv�Hj^
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���w�Hj[
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��{�Hh�)��}�(h�Kh�Kh�}��|�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��|�Hj�
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���{�Hj
  sh�Kh�hRh�h�)��}�(h�}��P{�Hj�
  sh�Kh�hRh�Nj0  h�)��}�(h�}��z�Hj�
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P{�Hj�
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj�
  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�
  sh�Kh�hRh�h�)��}�(h�}���Hj�
  sh�Kh�hRh�Nj0  h�)��}�(h�}���}�Hj�
  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���Hj�
  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj   sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�
  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�
  sh�Kh�hRh�h�)��}�(h�}���Hj  sh�Kh�hRh�Nj0  h�)��}�(h�}����Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���Hj  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj?  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj<  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj<  sh�Kh�hRh�h�)��}�(h�}���HjW  sh�Kh�hRh�Nj0  h�)��}�(h�}����HjZ  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���HjW  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�(�Hh�)��}�(h�Kh�Kh�}��P(�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P(�Hj~  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj{  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��(�Hj{  sh�Kh�hRh�h�)��}�(h�}��P%�Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}��%�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��P%�Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��+�Hh�)��}�(h�Kh�Kh�}��,�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��,�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���+�Hj�  sh�Kh�hRh�h�)��}�(h�}��P+�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��*�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P+�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��/�Hh�)��}�(h�Kh�Kh�}���/�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���/�Hj  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���/�Hj  sh�Kh�hRh�h�)��}�(h�}��/�Hj   sh�Kh�hRh�Nj0  h�)��}�(h�}���-�Hj#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}��/�Hj   sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P3�Hh�)��}�(h�Kh�Kh�}���Y�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���Y�HjG  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjD  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P3�HjD  sh�Kh�hRh�h�)��}�(h�}���2�Hje  sh�K h�hRh�Nj0  h�)��}�(h�}���1�Hjh  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���2�Hje  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PO�Hh�)��}�(h�Kh�Kh�}������Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}������Hj�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PO�Hj�  sh�Kh�hRh�h�)��}�(h�}���Pg�Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}��Z�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���Pg�Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�����Hh�)��}�(h�Kh�Kh�}��Ah�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Ah�Hj�  sh�Kh�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  Nubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}������Hj�  sh�Kh�hRh�h�)��}�(h�}���+��Hj�  sh�Kh�hRh�Nj0  h�)��}�(h�}��PW�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�Nubh�h�)��}�(h�}���+��Hj�  sh�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��Y�Hh�)��}�(h�Kh�Kh�}���X�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���X�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���Y�Hj  sh�Kh�hRh�h�)��}�(h�}��Y�Hj.  sh�K h�hRh�Nj0  h�)��}�(h�}��Pi�Hj1  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Y�Hj.  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�N�Hh�)��}�(h�Kh�Kh�}��PL�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PL�Hj[  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjX  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��N�HjX  sh�Kh�hRh�h�)��}�(h�}���G�Hjy  sh�K h�hRh�Nj0  h�)��}�(h�}��m�Hj|  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���G�Hjy  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��e�Hh�)��}�(h�Kh�Kh�}��F�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��F�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���e�Hj�  sh�Kh�hRh�h�)��}�(h�}��h�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���y�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��h�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Ў��Hh�)��}�(h�Kh�Kh�}������Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}������Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Ў��Hj�  sh�Kh�hRh�h�)��}�(h�}�����Hj  sh�K h�hRh�Nj0  h�)��}�(h�}���=��Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�
�Hh�)��}�(h�Kh�Kh�}��P�
�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�
�Hj<  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj9  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�
�Hj9  sh�Kh�hRh�h�)��}�(h�}����
�HjZ  sh�K h�hRh�Nj0  h�)��}�(h�}����
�Hj]  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����
�HjZ  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���
�Hh�)��}�(h�Kh�Kh�}����
�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����
�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����
�Hj�  sh�Kh�hRh�h�)��}�(h�}����
�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���
�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����
�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��
�Hh�)��}�(h�Kh�Kh�}����
�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����
�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���
�Hj�  sh�Kh�hRh�h�)��}�(h�}���
�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����
�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���
�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�
�Hh�)��}�(h�Kh�Kh�}����
�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����
�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�
�Hj  sh�Kh�hRh�h�)��}�(h�}��P�
�Hj;  sh�K h�hRh�Nj0  h�)��}�(h�}����
�Hj>  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�
�Hj;  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���
�Hh�)��}�(h�Kh�Kh�}����
�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����
�Hjh  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIje  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����
�Hje  sh�Kh�hRh�h�)��}�(h�}����
�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��P�
�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����
�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��(i�Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���(i�Hj�  sh�Kh�hRh�h�)��}�(h�}��i�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����
�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��i�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����Hj�  sh�Kh�hRh�h�)��}�(h�}��P��Hj  sh�K h�hRh�Nj0  h�)��}�(h�}��P��Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P��Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����Hh�)��}�(h�Kh�Kh�}�����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����HjI  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjF  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����HjF  sh�Kh�hRh�h�)��}�(h�}��P��Hjg  sh�K h�hRh�Nj0  h�)��}�(h�}�����Hjj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P��Hjg  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}�����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}�����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�  sh�Kh�hRh�h�)��}�(h�}����Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��#d�Hh�)��}�(h�Kh�Kh�}��P%d�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P%d�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���#d�Hj�  sh�Kh�hRh�h�)��}�(h�}�����Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}���l`�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���l`�Hj*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj'  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��Hj'  sh�Kh�hRh�h�)��}�(h�}�����HjH  sh�K h�hRh�Nj0  h�)��}�(h�}�����HjK  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����HjH  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���	�Hh�)��}�(h�Kh�Kh�}��P�	�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�	�Hju  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjr  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����	�Hjr  sh�Kh�hRh�h�)��}�(h�}��P�	�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���	�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�	�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��	�Hh�)��}�(h�Kh�Kh�}��P�	�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�	�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���	�Hj�  sh�Kh�hRh�h�)��}�(h�}��Ѕ	�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���	�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Ѕ	�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�	�Hh�)��}�(h�Kh�Kh�}���	�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���	�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�	�Hj  sh�Kh�hRh�h�)��}�(h�}���	�Hj)  sh�K h�hRh�Nj0  h�)��}�(h�}��Ї	�Hj,  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���	�Hj)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�	�Hh�)��}�(h�Kh�Kh�}��P�	�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�	�HjV  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjS  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�	�HjS  sh�Kh�hRh�h�)��}�(h�}��P�	�Hjt  sh�K h�hRh�Nj0  h�)��}�(h�}��P�	�Hjw  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�	�Hjt  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��	�Hh�)��}�(h�Kh�Kh�}��P�	�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�	�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���	�Hj�  sh�Kh�hRh�h�)��}�(h�}��P�	�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����	�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�	�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pa�Hh�)��}�(h�Kh�Kh�}��y�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��y�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�b�      j�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pa�Hj�  sh�Kh�hRh�h�)��}�(h�}��L�Hj
  sh�K h�hRh�Nj0  h�)��}�(h�}��P�	�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��L�Hj
  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��	�Hh�)��}�(h�Kh�Kh�}��5�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��5�Hj7  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj4  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���	�Hj4  sh�Kh�hRh�h�)��}�(h�}��P8�HjU  sh�K h�hRh�Nj0  h�)��}�(h�}��� �HjX  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P8�HjU  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�О�Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��О�Hj  sh�Kh�hRh�h�)��}�(h�}��С�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}�����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��С�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P^�Hh�)��}�(h�Kh�Kh�}��P�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P^�Hj�  sh�Kh�hRh�h�)��}�(h�}��PE�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���~�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PE�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��L�Hh�)��}�(h�Kh�Kh�}��PZ�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PZ�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���L�Hj  sh�Kh�hRh�h�)��}�(h�}��`�Hj6  sh�K h�hRh�Nj0  h�)��}�(h�}���O�Hj9  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��`�Hj6  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��X�Hh�)��}�(h�Kh�Kh�}���x�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���x�Hjc  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj`  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���X�Hj`  sh�Kh�hRh�h�)��}�(h�}���Z�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���v�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���Z�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PX�Hh�)��}�(h�Kh�Kh�}���i�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���i�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PX�Hj�  sh�Kh�hRh�h�)��}�(h�}��_�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��Ps�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��_�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��l�Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���l�Hj�  sh�Kh�hRh�h�)��}�(h�}���e�Hj  sh�K h�hRh�Nj0  h�)��}�(h�}���g�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���e�Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P*��Hh�)��}�(h�Kh�Kh�}��Ўe�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Ўe�HjD  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjA  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P*��HjA  sh�Kh�hRh�h�)��}�(h�}��=��Hjb  sh�K h�hRh�Nj0  h�)��}�(h�}��P9��Hje  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��=��Hjb  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��Hj�  sh�Kh�hRh�h�)��}�(h�}��P��Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��ŋ�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P��Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub����Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}�����Hj�  sh�Kh�hRh�h�)��}�(h�}����Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}��P7�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P7�Hj%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj"  sh�Kh�hRh�h�)��}�(h�}����HjC  sh�K h�hRh�Nj0  h�)��}�(h�}�����HjF  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����HjC  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Џ��Hh�)��}�(h�Kh�Kh�}��Е��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Е��Hjp  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjm  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Џ��Hjm  sh�Kh�hRh�h�)��}�(h�}��P���Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P���Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}��P��Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P��Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��Hj�  sh�Kh�hRh�h�)��}�(h�}�����Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}�����Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P��Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P��Hj  sh�Kh�hRh�h�)��}�(h�}��е�Hj$  sh�K h�hRh�Nj0  h�)��}�(h�}��P��Hj'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��е�Hj$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�\��Hh�)��}�(h�Kh�Kh�}���C�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���C�HjQ  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjN  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��\��HjN  sh�Kh�hRh�h�)��}�(h�}��A�Hjo  sh�K h�hRh�Nj0  h�)��}�(h�}��K��Hjr  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��A�Hjo  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�#�Hh�)��}�(h�Kh�Kh�}���Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��#�Hj�  sh�Kh�hRh�h�)��}�(h�}��P�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�4�Hh�)��}�(h�Kh�Kh�}���8�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���8�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��4�Hj�  sh�Kh�hRh�h�)��}�(h�}��P7�Hj  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P7�Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��9�Hh�)��}�(h�Kh�Kh�}���?�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���?�Hj2  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj/  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���9�Hj/  sh�Kh�hRh�h�)��}�(h�}��?�HjP  sh�K h�hRh�Nj0  h�)��}�(h�}��P9�HjS  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��?�HjP  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�B�Hh�)��}�(h�Kh�Kh�}���F�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���F�Hj}  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjz  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��B�Hjz  sh�Kh�hRh�h�)��}�(h�}��PE�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���@�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PE�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�H�Hh�)��}�(h�Kh�Kh�}��M�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��M�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��H�Hj�  sh�Kh�hRh�h�)��}�(h�}���L�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���I�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���L�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��N�Hh�)��}�(h�Kh�Kh�}���S�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���S�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���N�Hj  sh�Kh�hRh�h�)��}�(h�}��PS�Hj1  sh�K h�hRh�Nj0  h�)��}�(h�}��PP�Hj4  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PS�Hj1  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PT�Hh�)��}�(h�Kh�Kh�}���Y�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���Y�Hj^  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj[  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PT�Hj[  sh�Kh�hRh�h�)��}�(h�}���Y�Hj|  sh�K h�hRh�Nj0  h�)��}�(h�}��T�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���Y�Hj|  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��`�Hh�)��}�(h�Kh�Kh�}���[�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���[�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���`�Hj�  sh�Kh�hRh�h�)��}�(h�}���^�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��PZ�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���^�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��b�Hh�)��}�(h�Kh�Kh�}���g�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���g�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���b�Hj�  sh�Kh�hRh�h�)��}�(h�}��g�Hj  sh�K h�hRh�Nj0  h�)��}�(h�}��a�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��g�Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pi�Hh�)��}�(h�Kh�Kh�}��n�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��n�Hj?  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj<  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pi�Hj<  sh�Kh�hRh�h�)��}�(h�}���l�Hj]  sh�K h�hRh�Nj0  h�)��}�(h�}���j�Hj`  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���l�Hj]  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pp�Hh�)��}�(h�Kh�Kh�}���t�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���t�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pp�Hj�  sh�Kh�hRh�h�)��}�(h�}���s�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���n�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���s�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��v�Hh�)��}�(h�Kh�Kh�}���{�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���{�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���v�Hj�  sh�Kh�hRh�h�)��}�(h�}��P{�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��Pu�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P{�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��Hh�)��}�(h�Kh�Kh�}���Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���Hj   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���Hj  sh�Kh�hRh�h�)��}�(h�}����Hj>  sh�K h�hRh�Nj0  h�)��}�(h�}���|�HjA  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj>  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�Hh�)��}�(h�Kh�Kh�}��P
�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P
�Hjk  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjh  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�Hjh  sh�Kh�hRh�h�)��}�(h�}���	�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���	�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��"�Hh�)��}�(h�Kh�Kh�}��#�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��#�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���"�Hj�  sh�Kh�hRh�h�)��}�(h�}���"�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���"�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��'�Hh�)��}�(h�Kh�Kh�}��(�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��(�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���'�Hj�  sh�Kh�hRh�h�)��}�(h�}���'�Hj  sh�K h�hRh�Nj0  h�)��}�(h�}���&�Hj"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���'�Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�*�Hh�)��}�(h�Kh�Kh�}���.�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���.�HjL  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjI  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��*�HjI  sh�Kh�hRh�h�)��}�(h�}��.�Hjj  sh�K h�hRh�Nj0  h�)��}�(h�}���(�Hjm  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��.�Hjj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P2�Hh�)��}�(h�Kh�Kh�}���5�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���5�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P2�Hj�  sh�Kh�hRh�h�)��}�(h�}��P4�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���4�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P4�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��9�Hh�)��}�(h�Kh�Kh�}��=�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��=�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���9�Hj�  sh�Kh�hRh�h�)��}�(h�}���<�Hj   sh�K h�hRh�Nj0  h�)��}�(h�}���:�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���<�Hj   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�A�Hh�)��}�(h�Kh�Kh�}��PD�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PD�Hj-  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj*  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��A�Hj*  sh�Kh�hRh�h�)��}�(h�}��C�HjK  sh�K h�hRh�Nj0  h�)��}�(h�}���@�HjN  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��C�HjK  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�F�Hh�)��}�(h�Kh�Kh�}���J�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���J�Hjx  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIju  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��F�Hju  sh�Kh�hRh�h�)��}�(h�}���I�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���G�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���I�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��K�Hh�)��}�(h�Kh�Kh�}��PQ�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PQ�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���K�Hj�  sh�Kh�hRh�h�)��}�(h�}��Q�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��PN�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Q�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�R�Hh�)��}�(h�Kh�Kh�}��PV�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PV�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��R�Hj  sh�Kh�hRh�h�)��}�(h�}��PU�Hj,  sh�K h�hRh�Nj0  h�)��}�(h�}���R�Hj/  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PU�Hj,  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Z�Hh�)��}�(h�Kh�Kh�}��\�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��\�HjY  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjV  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Z�HjV  sh�Kh�hRh�h�)��}�(h�}��[�Hjw  sh�K h�hRh�Nj0  h�)��}�(h�}���W�Hjz  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��[�Hjw  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��^�Hh�)��}�(h�Kh�Kh�}���c�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���c�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���^�Hj�  sh�Kh�hRh�h�)��}�(h�}��Pb�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}��P`�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Pb�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��e�Hh�)��}�(h�Kh�Kh�}���j�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���j�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���e�Hj�  sh�Kh�hRh�h�)��}�(h�}��Pj�Hj  sh�K h�hRh�Nj0  h�)��}�(h�}��g�Hj  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Pj�Hj  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��k�Hh�)��}�(h�Kh�Kh�}��Pq�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pq�Hj:  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj7  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���k�Hj7  sh�Kh�hRh�h�)��}�(h�}��q�HjX  sh�K h�hRh�Nj0  h�)��}�(h�}��Pn�Hj[  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��q�HjX  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Ps�Hh�)��}�(h�Kh�Kh�}��Px�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Px�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Ps�Hj�  sh�Kh�hRh�h�)��}�(h�}��x�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���q�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��x�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�z�Hh�)��}�(h�Kh�Kh�}���~�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���~�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��z�Hj�  sh�Kh�hRh�h�)��}�(h�}���}�Hj�  sh�K h�hRh�Nj0  h�)��}�(h�}���{�Hj�  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���}�Hj�  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��B�Hh�)��}�(h�Kh�Kh�}��PF�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PF�Hj   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���B�Hj   sh�Kh�hRh�h�)��}�(h�}���E�Hj9   sh�K h�hRh�Nj0  h�)��}�(h�}��P@�Hj<   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���E�Hj9   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��G�Hh�)��}�(h�Kh�Kh�}��M�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��M�Hjf   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjc   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���G�Hjc   sh�Kh�hRh�h�)��}�(h�}���L�Hj�   sh�K h�hRh�Nj0  h�)��}�(h�}��E�Hj�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���L�Hj�   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��O�Hh�)��}�(h�Kh�Kh�}���S�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���S�Hj�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���O�Hj�   sh�Kh�hRh�h�)��}�(h�}��PR�Hj�   sh�K h�hRh�Nj0  h�)��}�(h�}���L�Hj�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PR�Hj�   sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��V�Hh�)��}�(h�Kh�Kh�}���X�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���X�Hj�   sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�   j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���V�Hj�   sh�Kh�hRh�h�)��}�(h�}���W�Hj!  sh�K h�hRh�Nj0  h�)��}�(h�}��PS�Hj!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���W�Hj!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P[�Hh�)��}�(h�Kh�Kh�}���_�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���_�HjG!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjD!  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P[�HjD!  sh�Kh�hRh�h�)��}�(h�}���^�Hje!  sh�K h�hRh�Nj0  h�)��}�(h�}���Y�Hjh!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���^�Hje!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pa�Hh�)��}�(h�Kh�Kh�}��f�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��f�Hj�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�!  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pa�Hj�!  sh�Kh�hRh�h�)��}�(h�}���d�Hj�!  sh�K h�hRh�Nj0  h�)��}�(h�}���b�Hj�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���d�Hj�!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��f�Hh�)��}�(h�Kh�Kh�}��Pl�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pl�Hj�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�!  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���f�Hj�!  sh�Kh�hRh�h�)��}�(h�}��k�Hj�!  sh�K h�hRh�Nj0  h�)��}�(h�}���e�Hj�!  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��k�Hj�!  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�l�Hh�)��}�(h�Kh�Kh�}��Pr�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pr�Hj("  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj%"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��l�Hj%"  sh�Kh�hRh�h�)��}�(h�}��r�HjF"  sh�K h�hRh�Nj0  h�)��}�(h�}��Po�HjI"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��r�HjF"  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Pt�Hh�)��}�(h�Kh�Kh�}��y�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��y�Hjs"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjp"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Pt�Hjp"  sh�Kh�hRh�h�)��}�(h�}���w�Hj�"  sh�K h�hRh�Nj0  h�)��}�(h�}���u�Hj�"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���w�Hj�"  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P|�Hh�)��}�(h�Kh�Kh�}��P�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�Hj�"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�"  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P|�Hj�"  sh�Kh�hRh�h�)��}�(h�}���Hj�"  sh�K h�hRh�Nj0  h�)��}�(h�}��Ps�Hj�"  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���Hj�"  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��B�Hh�)��}�(h�Kh�Kh�}���E�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���E�Hj	#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���B�Hj#  sh�Kh�hRh�h�)��}�(h�}���D�Hj'#  sh�K h�hRh�Nj0  h�)��}�(h�}��P@�Hj*#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���D�Hj'#  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PF�Hh�)��}�(h�Kh�Kh�}��L�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��L�HjT#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjQ#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PF�HjQ#  sh�Kh�hRh�h�)��}�(h�}���J�Hjr#  sh�K h�hRh�Nj0  h�)��}�(h�}��E�Hju#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���J�Hjr#  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PO�Hh�)��}�(h�Kh�Kh�}��PQ�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��PQ�Hj�#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PO�Hj�#  sh�Kh�hRh�h�)��}�(h�}��PP�Hj�#  sh�K h�hRh�Nj0  h�)��}�(h�}���K�Hj�#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PP�Hj�#  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�U�Hh�)��}�(h�Kh�Kh�}���X�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���X�Hj�#  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�#  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��U�Hj�#  sh�Kh�hRh�h�)��}�(h�}��PX�Hj$  sh�K h�hRh�Nj0  h�)��}�(h�}���R�Hj$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PX�Hj$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PZ�Hh�)��}�(h�Kh�Kh�}��_�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��_�Hj5$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj2$  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PZ�Hj2$  sh�Kh�hRh�h�)��}�(h�}���]�HjS$  sh�K h�hRh�Nj0  h�)��}�(h�}���[�HjV$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���]�HjS$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�a�Hh�)��}�(h�Kh�Kh�}���e�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���e�Hj�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj}$  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��a�Hj}$  sh�Kh�hRh�h�)��}�(h�}��Pd�Hj�$  sh�K h�hRh�Nj0  h�)��}�(h�}���_�Hj�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Pd�Hj�$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�f�Hh�)��}�(h�Kh�Kh�}���k�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���k�Hj�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�$  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��f�Hj�$  sh�Kh�hRh�h�)��}�(h�}���k�Hj�$  sh�K h�hRh�Nj0  h�)��}�(h�}���h�Hj�$  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���k�Hj�$  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��l�Hh�)��}�(h�Kh�Kh�}��Pr�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��Pr�Hj%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���l�Hj%  sh�Kh�hRh�h�)��}�(h�}��r�Hj4%  sh�K h�hRh�Nj0  h�)��}�(h�}��Po�Hj7%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��r�Hj4%  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�t�Hh�)��}�(h�Kh�Kh�}���x�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���x�Hja%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj^%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��t�Hj^%  sh�Kh�hRh�h�)��}�(h�}���w�Hj%  sh�K h�hRh�Nj0  h�)��}�(h�}���u�Hj�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���w�Hj%  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Py�Hh�)��}�(h�Kh�Kh�}���Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���Hj�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Py�Hj�%  sh�Kh�hRh�h�)��}�(h�}���~�Hj�%  sh�K h�hRh�Nj0  h�)��}�(h�}��|�Hj�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���~�Hj�%  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P �Hh�)��}�(h�Kh�Kh�}��P�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�Hj�%  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�%  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P �Hj�%  sh�Kh�hRh�h�)��}�(h�}����Hj&  sh�K h�hRh�Nj0  h�)��}�(h�}��� �Hj&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����HjB&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj?&  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj?&  sh�Kh�hRh�h�)��}�(h�}��P�Hj`&  sh�K h�hRh�Nj0  h�)��}�(h�}���	�Hjc&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�Hj`&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}��P�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��P�Hj�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�&  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj�&  sh�Kh�hRh�h�)��}�(h�}����Hj�&  sh�K h�hRh�Nj0  h�)��}�(h�}���Hj�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj�&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�&  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubs�      h�Kh�hRh�h�)��}�(h�Kh�Kh�}���Hj�&  sh�Kh�hRh�h�)��}�(h�}��P�Hj�&  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj�&  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P�Hj�&  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub���Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj#'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj '  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}����Hj '  sh�Kh�hRh�h�)��}�(h�}����HjA'  sh�K h�hRh�Nj0  h�)��}�(h�}���HjD'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����HjA'  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P!�Hh�)��}�(h�Kh�Kh�}��&�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��&�Hjn'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjk'  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P!�Hjk'  sh�Kh�hRh�h�)��}�(h�}���$�Hj�'  sh�K h�hRh�Nj0  h�)��}�(h�}���"�Hj�'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���$�Hj�'  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��%�Hh�)��}�(h�Kh�Kh�}���,�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���,�Hj�'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�'  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���%�Hj�'  sh�Kh�hRh�h�)��}�(h�}��,�Hj�'  sh�K h�hRh�Nj0  h�)��}�(h�}��)�Hj�'  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��,�Hj�'  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��.�Hh�)��}�(h�Kh�Kh�}���3�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���3�Hj(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���.�Hj(  sh�Kh�hRh�h�)��}�(h�}��P3�Hj"(  sh�K h�hRh�Nj0  h�)��}�(h�}��-�Hj%(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��P3�Hj"(  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�7�Hh�)��}�(h�Kh�Kh�}��9�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}��9�HjO(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjL(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��7�HjL(  sh�Kh�hRh�h�)��}�(h�}��8�Hjm(  sh�K h�hRh�Nj0  h�)��}�(h�}���3�Hjp(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��8�Hjm(  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��9�Hh�)��}�(h�Kh�Kh�}���?�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���?�Hj�(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���9�Hj�(  sh�Kh�hRh�h�)��}�(h�}���>�Hj�(  sh�K h�hRh�Nj0  h�)��}�(h�}��=�Hj�(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���>�Hj�(  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��@�Hh�)��}�(h�Kh�Kh�}���F�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���F�Hj�(  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�(  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���@�Hj�(  sh�Kh�hRh�h�)��}�(h�}��PF�Hj)  sh�K h�hRh�Nj0  h�)��}�(h�}���C�Hj)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PF�Hj)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��E�Hh�)��}�(h�Kh�Kh�}���L�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���L�Hj0)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj-)  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���E�Hj-)  sh�Kh�hRh�h�)��}�(h�}��PL�HjN)  sh�K h�hRh�Nj0  h�)��}�(h�}���I�HjQ)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��PL�HjN)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�PO�Hh�)��}�(h�Kh�Kh�}���R�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���R�Hj{)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjx)  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��PO�Hjx)  sh�Kh�hRh�h�)��}�(h�}���R�Hj�)  sh�K h�hRh�Nj0  h�)��}�(h�}���K�Hj�)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���R�Hj�)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub��S�Hh�)��}�(h�Kh�Kh�}���Y�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���Y�Hj�)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj�)  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}���S�Hj�)  sh�Kh�hRh�h�)��}�(h�}��Y�Hj�)  sh�K h�hRh�Nj0  h�)��}�(h�}��W�Hj�)  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}��Y�Hj�)  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�Z�Hh�)��}�(h�Kh�Kh�}���^�Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}���^�Hj*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIj*  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��Z�Hj*  sh�Kh�hRh�h�)��}�(h�}���]�Hj/*  sh�K h�hRh�Nj0  h�)��}�(h�}���\�Hj2*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}���]�Hj/*  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ub�P�Hh�)��}�(h�Kh�Kh�}����Hh�)��}�(h�}�h�Kh�hRj�  h�)��}�(h�}����Hj\*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubhIjY*  j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�Kh�hRh�h�)��}�(h�Kh�Kh�}��P�HjY*  sh�Kh�hRh�h�)��}�(h�}����Hjz*  sh�K h�hRh�Nj0  h�)��}�(h�}����Hj}*  sh�K h�hRj�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hjz*  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bububh�h�ubuh�Kh�hRh�Nj0  h�h�hhK ��h��R�(KKK��h!�CH      Y@        �8��8V�@             xz@9��8��I@                      �?�t�bubsh�Kh�hRj�  h�hIh�j�  hhK ��h��R�(KKK��h!�C �8��8V�@9��8��I@�8��8v�@�q�q�}@�t�bubsh�K h�hRj�  hhK ��h��R�(KKK��h!�C �������?(\���(�?�������?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bub�_originalPosition�h�)��}�(h�}�h�Kh�hRj�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bub�_aspect�h7�_adjustable��box��_anchor��C��_stale_viewlims�}�(h~�h��u�_sharex�N�_sharey�h>�bbox�h��dataLim�h�)��}�(h�}�h�Kh�hRj�  hhK ��h��R�(KKK��h!�C         ���`C!�     �E@ڜ��H��?�t�bj�  hhK ��h��R�(KK��h!�C      �?�>���q?�t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �      �      ��      ���t�bub�_viewLim�j	  �
transScale�j�  �	transAxes�h��transLimits�j	  �	transData�h��_xaxis_transform�h��_yaxis_transform�j	  �_subplotspec�N�_box_aspect�N�_axes_locator��	functools��partial���h��$mpl_toolkits.axes_grid1.axes_divider��AxesDivider���)��}�(hBh>�_xref��!mpl_toolkits.axes_grid1.axes_size��AxesX���)��}�(hBh>j�*  G?�      �_ref_ax�Nub�_yref�j+  �AxesY���)��}�(hBh>j�*  G?�      j+  Nub�_fig�hG�_pos�N�_horizontal�]�(j+  j+  �Fixed���)��}��
fixed_size�G?�������sbj+  )��}�j+  Ksbe�	_vertical�]�j+  aj�*  j�*  j�*  N�
_xrefindex�K �
_yrefindex�K �_locator�Nub�_locate���R���R�(j(+  (KK KKt�}�}��get_subplotspec�h�j+  j.+  ��R�st�b�	_children�]�(�matplotlib.patches��	Rectangle���)��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQ�
_nolegend_�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx��_hatch_color�(G        G        G        G?�      t��_fill���_original_edgecolor�N�
_edgecolor�(G        G        G        G        t��_original_facecolor�hhK ��h��R�(KK��h!�C �?�������?TTTTTT�?      �?�t�b�
_facecolor�(G?�G?ܜ�����G?�TTTTTTG?�      t��
_linewidth�G?�333333�_unscaled_dash_pattern�K N���_dash_pattern�G        N���
_linestyle��solid��_antialiased���_hatch�N�	_capstyle��matplotlib._enums��CapStyle����butt���R��
_joinstyle�jb+  �	JoinStyle����miter���R��_x0�jE+  �_y0�h0h!C���`C!⿔��R��_width�h0h!C       @���R��_height�h0h!C@����[�?���R��angle�G        �_rotation_point��xy��_aspect_ratio_correction�G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj[  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�+  jo+  h0h!Cr��id^῔��R�js+  h0h!C        ���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�+  jo+  h0h!C�iLr��࿔��R�js+  h0h!C      �?���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�+  jo+  h0h!C�H0�L�߿���R�js+  h0h!C        ���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj<  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�+  jo+  h0h!C	���+޿���R�js+  h0h!C      �?���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j ,  jo+  h0h!C3_ѥܿ���R�js+  h0h!C       @���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j,  jo+  h0h!C$��* ۿ���R�js+  h0h!C      @���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j:,  jo+  h0h!C0�<U�ٿ���R�js+  h0h!C      @���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjh  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jW,  jo+  h0h!C;�%N�ؿ���R�js+  h0h!C      @���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jt,  jo+  h0h!CI�_ֿَ���R�js+  h0h!C        ���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�,  jo+  h0h!CV|Tq	տ���R�js+  h0h!C       @���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjI  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�,  jo+  h0h!Ca��]�ӿ���R�js+  h0h!C      @���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�,  jo+  h0h!Cof����ѿ���R�js+  h0h!C      @���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�,  jo+  h0h!Cz���wп���R�js+  h0h!C      *@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj*  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j-  jo+  h0h!C�doG�Ϳ���R�js+  h0h!C      &@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNju  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j"-  jo+  h0h!C'�����ʿ���R�js+  h0h!C       @���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j?-  jo+  h0h!CAuµO�ǿ���R�js+  h0h!C      &@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j\-  jo+  h0h!C\_����Ŀ���R�js+  h0h!C      3@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjV  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jy-  jo+  h0h!CsI �W������R�js+  h0h!C      4@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�-  jo+  h0h!Cg�>�U�����R�js+  h0h!C      >@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�-  jo+  h0h!CJ;���>�����R�js+  h0h!C      :@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj7  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�-  jo+  h0h!C�Z��'�����R�js+  h0h!C      ?@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�-  jo+  h0h!C`�o#�!�����R�js+  h0h!C      E@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j
.  jo+  h0h!C��V`e瓿���R�js+  h0h!C     �E@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j'.  jo+  h0h!C�>���q?���R�js+  h0h!C      >@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjc  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jD.  jo+  h0h!C�~�lXМ?���R�js+  h0h!C      <@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  ja.  jo+  h0h!C�����?���R�js+  h0h!C      4@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j~.  jo+  h0h!CP�r�b�?���R�js+  h0h!C      6@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjD  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�.  jo+  h0h!C #H�x�?���R�js+  h0h!C      =@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�.  jo+  h0h!C�N����?���R�js+  h0h!C      5@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�.  jo+  h0h!C`��]v��?���R�js+  h0h!C      2@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj%  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�.  jo+  h0h!CD�}:���?���R�js+  h0h!C      1@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjp  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j/  jo+  h0h!C,�Nn��?���R�js+  h0h!C      ,@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j,/  jo+  h0h!C�����?���R�js+  h0h!C      (@���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jI/  jo+  h0h!C���e�?���R�js+  h0h!C      *@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjQ  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jf/  jo+  h0h!Cp��p�?���R�js+  h0h!C        ���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�/  jo+  h0h!Cd�I�.��?���R�js+  h0h!C      &@���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�/  jo+  h0h!CX+����?���R�js+  h0h!C      �?���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj2  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�/  jo+  h0h!CJ�����?���R�js+  h0h!C      @���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj}  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�/  jo+  h0h!C>A��h�?���R�js+  h0h!C      �?���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�/  jo+  h0h!C2��~&��?���R�js+  h0h!C       @���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j0  jo+  h0h!C$WTm�(�?���R�js+  h0h!C      �?���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj^  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j10  jo+  h0h!C�[���?���R�js+  h0h!C       @���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jN0  jo+  h0h!Cm%J`4�?���R�js+  h0h!C      �?���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jk0  jo+  h0h!C ��8��?���R�js+  h0h!C        ���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj?  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�0  jo+  h0h!CzA{��?���R�js+  h0h!C        ���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�0  jo+  h0h!C�
���?���R�js+  h0h!C      �?���R�jw+  h0h!C ����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�0  jo+  h0h!Cl�����?���R�js+  h0h!C        ���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj   hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�0  jo+  h0h!C���h�?���R�js+  h0h!C      �?���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjk  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  jR+  jV+  (G?�G?ܜ�����G?�TTTTTTG?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�0  jo+  h0h!C`WL�i+�?���R�js+  h0h!C      �?���R�jw+  h0h!C@����[�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  hhK ��h��R�(KK��h!�C �������?xxxxxx�?�������?      �?�t�bjV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j1  jo+  h0h!C(�R�J߿���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j<1  jo+  h0h!COajJ��ݿ���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjL  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jY1  jo+  h0h!Ctځ���ܿ���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jv1  jo+  h0h!C�S�A]ۿ���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�1  jo+  h0h!C�̰|�%ڿ���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj-  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�1  jo+  h0h!C�E���ؿ���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjx  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�1  jo+  h0h!C��H7�׿���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�1  jo+  h0h!C68���ֿ���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j2  jo+  h0h!C\��Hտ���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjY  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j$2  jo+  h0h!C�*&{-Կ���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jA2  jo+  h0h!C��=���ҿ���R�js+  h0h!C       @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j^2  jo+  h0h!C�UG|�ѿ���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj:  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j{2  jo+  h0h!C��l�#kп���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�2  jo+  h0h!C<'�gο���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�2  jo+  h0h!C�7���˿���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj   hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�2  jo+  h0h!C�f�3�ɿ���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjf   hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�2  jo+  h0h!C"����ǿ���R�js+  h0h!C       @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�   hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j3  jo+  h0h!Cp��WѬĿ���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�   hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j)3  jo+  h0h!C���# >¿���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjG!  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jF3  jo+  h0h!C�C�ݞ�����R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�!  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jc3  jo+  h0h!C�|�x{������R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�!  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�3  jo+  h0h!CHa�䵿���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj("  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�3  jo+  h0h!C�E]�������R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjs"  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�3  jo+  h0h!C�Tv��R�����R�js+  h0h!C       @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�"  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�3  jo+  h0h!C`<dh�/�����R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj	#  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�3  jo+  h0h!C����{t�����R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjT#  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j4  jo+  h0h!C�=Y��v�?���R�js+  h0h!C      $@���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�#  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j.4  jo+  h0h!C`5s�0�?���R�js+  h0h!C       @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�#  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jK4  jo+  h0h!C �ވ/S�?���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj5$  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jh4  jo+  h0h!C�y,��?���R�js+  h0h!C       @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�$  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�4  jo+  h0h!CP���\�?���R�js+  h0h!C       @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�$  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�4  jo+  h0h!C��U����?���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj%  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�4  jo+  h0h!C��b!��?���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNja%  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�4  jo+  h0h!C��L�A>�?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�%  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�4  jo+  h0h!Cp��?���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�%  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j5  jo+  h0h!C$�L��?���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjB&  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j35  jo+  h0h!C���U��?���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�&  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jP5  jo+  h0h!C�*����?���R�js+  h0h!C      @���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�&  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jm5  jo+  h0h!C<8b�g�?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj#'  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�5  jo+  h0h!C���4k�?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjn'  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�5  jo+  h0h!C�)(���?���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�'  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�5  jo+  h0h!C�������?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj(  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�5  jo+  h0h!C�7�[>�?���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNjO(  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�5  jo+  h0h!C^����H�?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�(  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j6  jo+  h0h!C8E����?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�(  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j86  jo+  h0h!C̌)H��?���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj0)  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jU6  jo+  h0h!C�Ruà��?���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj{)  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  jr6  jo+  h0h!C��]]�%�?���R�js+  h0h!C        ���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj�)  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�6  jo+  h0h!C�`F�Q]�?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNj*  hONhP�hQj9+  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�h0h!C        ���R�a]�����hx�jI+  jJ+  jK+  �jL+  NjM+  jN+  jO+  j1  jV+  (G?�������G?�xxxxxxG?�������G?�      t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  j�6  jo+  h0h!Cv�.����?���R�js+  h0h!C      �?���R�jw+  h0h!C�m���u�?���R�j{+  G        j|+  j}+  j~+  G?�      ub�matplotlib.lines��Line2D���)��}�(h@�hANhBh�hChGhIj	  hJ�hK�hL�hMNhNj\*  hONhP�hQ�	_child100�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j3+  �remove���R�hjNhkNhlNhmNhnhohphs]�]�����hx��_dashcapstyle�jg+  �_dashjoinstyle�jj+  �round���R��_solidjoinstyle�j�6  �_solidcapstyle�jd+  j�6  ��R��_linestyles�N�
_drawstyle��default�jX+  G?�      jY+  K N��j[+  G        N��j]+  �-��	_invalidx���_color��#111111��_marker��matplotlib.markers��MarkerStyle���)��}�(�_marker_function�h�j�6  �_set_nothing���R��_user_transform�N�_user_capstyle�N�_user_joinstyle�N�
_fillstyle��full�j�6  �None�j#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�C �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nub�	_alt_path�N�_alt_transform�N�_snap_threshold�Njh+  j�6  ja+  jg+  �_filled��ub�	_gapcolor�N�
_markevery�N�_markersize�G@      j_+  ��_markeredgecolor��auto��_markeredgewidth�G        �_markerfacecolor��auto��_markerfacecoloralt��none��	_invalidy���_pickradius�K�
ind_offset�K �_xorig�]�(K Ke�_yorig�]�(K K ej�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�b�_xy�hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  j>  j5  j;  �	_subslice���	_x_filled�Nube�
_colorbars�]��spines��matplotlib.spines��Spines���)��}�(�left�j(7  �Spine���)��}�(h@�hANhBh�hChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  (G?陙����G?陙����G?陙����G?�      t�jK+  �jL+  �.8�jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jd+  �
projecting���R�jh+  jm+  �
spine_type�j-7  �axis��matplotlib.axis��YAxis���)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj?  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx��_remove_overlapping_locs���isDefault_label���major�jD7  �Ticker���)��}�(j%+  �matplotlib.ticker��AutoLocator���)��}�(�_nbins�h7�
_symmetric���_prune�N�_min_n_ticks�K�_steps�hhK ��h��R�(KK��h!�C(      �?       @      @      @      $@�t�b�_extended_steps�hhK ��h��R�(KK
��h!�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�b�_integer��jC7  jF7  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jR7  �jS7  �jT7  jW7  �minor�jV7  )��}�(j%+  jY7  �NullLocator���)��}�jC7  jq7  sb�
_formatter�jY7  �NullFormatter���)��}�(jC7  jq7  �locs�hhK ��h��R�(KK ��h!�j�6  t�bub�_locator_is_default���_formatter_is_default��ubhchZ)��}�(h]]��units�ah`hbhc}�j�7  }�K j+  h�h>�_unit_change_handler���R���R�(j�7  h���}��event��builtins��object���)��sNt�bssheKhfNhg��(K �ub�_autolabelpos���label��matplotlib.text��Text���)��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  h0h!C������7@���R�j�  G?�      �_text��	Residuals�j�6  �.15��_fontproperties��matplotlib.font_manager��FontProperties���)��}�(�_family�]��
sans-serif�a�_slant��normal��_variant��normal��_weight��normal��_stretch��normal��_file�N�_size�G@&      �_math_fontfamily��
dejavusans�ub�_usetex���_parse_math���_wrap���_verticalalignment��bottom��_horizontalalignment��center��_multialignment�N�	_rotation�G@V�     �_transform_rotates_text���_bbox_patch�N�	_renderer�N�_linespacing�G?�333333�_rotation_mode��anchor�j_+  �ub�
offsetText�j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  h0h!Cr�q�}@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  �      j�7  j�7  j�7  j�7  j�7  j�7  �normal�j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  �baseline�j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ub�labelpad�G@      j
7  K�_major_tick_kw�}�(�gridOn���tick1On���tick2On���label1On���label2On��u�_minor_tick_kw�}�(j�7  �j�7  �j�7  �j�7  �j�7  �u�	converter�Nj�7  N�_autoscale_on���label_position�j-7  �offset_text_position�j-7  �zorder�G?�      �_scale��matplotlib.scale��LinearScale���)���
majorTicks�]�(jD7  �YTick���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj#  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx��_loc�h0h!C������鿔��R��_major��j�7  G        js+  G?�      �	_base_pad�G@      �_labelrotation�j�6  K ���_zorder�G@ z�G��	tick1line�j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  �None�j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j,8  �_set_tickleft���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j8  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nub�	tick2line�j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jR8  �_set_tickright���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j8  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nub�gridline�j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�jp8  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j8  ��j	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nub�label1�j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j8  j�7  �−0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  �center_baseline�j�7  �right�j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ub�label2�j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j8  j�7  j�8  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ub�_tickdir��out��_pad�G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333㿔��R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�8  j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�8  ��j	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C433333㿔t�bj7  hhK ��h��R�(KKK��h!�C        433333㿔t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        433333㿔t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j9  jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�8  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j9  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�8  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�433333㿔t�bj7  hhK ��h��R�(KKK��h!�C         433333�      �?433333㿔t�bj#  j�  j5  j�  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�8  j�7  �−0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�8  j�7  jE9  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ٿ���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j)8  j[+  j*8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  jb9  ��j	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C        ������ٿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        ������ٿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jP8  j[+  jQ8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  jb9  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jn8  j[+  jo8  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  jb9  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ٿ������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ٿ      �?������ٿ�t�bj#  j
  j5  j  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  jb9  j�7  �−0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  jb9  j�7  j�9  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ɿ���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j)8  j[+  j*8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j:  ��j	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C        ������ɿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        ������ɿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jP8  j[+  jQ8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j:  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jn8  j[+  jo8  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j:  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ɿ������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ɿ      �?������ɿ�t�bj#  j  j5  j  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j:  j�7  �−0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j:  j�7  j�:  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C        ���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j)8  j[+  j*8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�:  ��j	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C                �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jP8  j[+  jQ8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�:  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jn8  j[+  jo8  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�:  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�bj7  hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  j(  j5  j%  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�:  j�7  �0.0�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�:  j�7  jm;  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j)8  j[+  j*8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�;  ��j	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C        �������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jP8  j[+  jQ8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�;  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jn8  j[+  jo8  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�;  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  j7  j5  j4  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�;  j�7  �0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�;  j�7  j%<  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j)8  j[+  j*8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  jB<  ��j	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C        �������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jP8  j[+  jQ8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  jB<  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jn8  j[+  jo8  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  jB<  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  jF  j5  jC  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  jB<  j�7  �0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  jB<  j�7  j�<  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333�?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j)8  j[+  j*8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�<  ��j	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C433333�?�t�bj7  hhK ��h��R�(KKK��h!�C        433333�?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        433333�?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jP8  j[+  jQ8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�<  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jn8  j[+  jo8  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�<  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�?433333�?�t�bj7  hhK ��h��R�(KKK��h!�C         433333�?      �?433333�?�t�bj#  jU  j5  jR  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�<  j�7  �0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�<  j�7  j�=  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j)8  j[+  j*8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�=  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jP8  j[+  jQ8  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�=  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjb  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jn8  j[+  jo8  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�=  ��j	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�=  j�7  �0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�=  j�7  j7>  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ube�
minorTicks�]�j8  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj7  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        js+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jb>  j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�K aj7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j~>  jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�Kaj7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMG?�      hNjv  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�>  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  ]�(K K ej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@333333ubaububj�7  jY7  �ScalarFormatter���)��}�(�_offset_threshold�K�offset�K �
_useOffset��j�7  ��_useMathText���orderOfMagnitude�K �format��%1.1f��_scientific���_powerlimits�]�(J����Ke�
_useLocale��jC7  jq7  j�7  hhK ��h��R�(KK	��h!�CH�������433333㿚�����ٿ������ɿ        �������?�������?433333�?�������?�t�bubj�7  �j�7  �ubj|7  j}7  hchZ)��}�(h]]�j�7  ah`hbhc}�j�7  }�K j+  h�h�j�7  ��R���R�(j�>  h���}�j�7  j�7  )��sNt�bssheKhfNhg��(K �ubj�7  �j�7  j�7  )��}�(h@�hANhBNhChGhIjk	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  h0h!C�q�)�@���R�j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@&      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G@V�     j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�7  j_+  �ubj�7  j�7  )��}�(h@�hANhBNhChGhIjw	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  h0h!Cr�q�}@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�7  G@      j
7  Kj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  Nj�7  Nj�7  �j�7  j-7  j�7  j-7  j�7  G?�      j 8  j8  j8  ]�(j8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj~  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������鿔��R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j5?  j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j&?  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jQ?  jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j&?  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�jm?  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j&?  ��j	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j&?  j�7  �−0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j&?  j�7  j�?  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333㿔��R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�?  j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�?  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�?  jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�?  ��j	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C433333㿔t�bj7  hhK ��h��R�(KKK��h!�C      �?433333㿔t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?433333㿔t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNjG  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j@  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�?  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�433333㿔t�bj7  hhK ��h��R�(KKK��h!�C         433333�      �?433333㿔t�bj#  jM  j5  jJ  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�?  j�7  �−0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�?  j�7  j;@  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ٿ���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j3?  j[+  j4?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  jX@  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jO?  j[+  jP?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  jX@  ��j	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C      �?������ٿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?������ٿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jk?  j[+  jl?  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  jX@  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ٿ������ٿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ٿ      �?������ٿ�t�bj#  j\  j5  jY  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  jX@  j�7  �−0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  jX@  j�7  j�@  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C������ɿ���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j3?  j[+  j4?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  jA  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jO?  j[+  jP?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  jA  ��j	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C      �?������ɿ�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?������ɿ�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jk?  j[+  jl?  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  jA  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C������ɿ������ɿ�t�bj7  hhK ��h��R�(KKK��h!�C         ������ɿ      �?������ɿ�t�bj#  jk  j5  jh  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  jA  j�7  �−0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  jA  j�7  j�A  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C        ���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j3?  j[+  j4?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�A  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jO?  j[+  jP?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�A  ��j	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jk?  j[+  jl?  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�A  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�bj7  hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  jz  j5  jw  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�A  j�7  �0.0�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�A  j�7  jcB  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j3?  j[+  j4?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�B  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jO?  j[+  jP?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�B  ��j	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jk?  j[+  jl?  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�B  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  j�  j5  j�  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�B  j�7  �0.2�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�B  j�7  jC  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j3?  j[+  j4?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j8C  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jO?  j[+  jP?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j8C  ��j	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�t�bj7  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?�������?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jk?  j[+  jl?  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j8C  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C�������?�������?�t�bj7  hhK ��h��R�(KKK��h!�C         �������?      �?�������?�t�bj#  j�  j5  j�  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j8C  j�7  �0.4�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j8C  j�7  j�C  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C433333�?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j3?  j[+  j4?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�C  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jO?  j[+  jP?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  �      G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�C  ��j	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C433333�?�t�bj7  hhK ��h��R�(KKK��h!�C      �?433333�?�t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?433333�?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jk?  j[+  jl?  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�C  ��j	7  �j�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C433333�?433333�?�t�bj7  hhK ��h��R�(KKK��h!�C         433333�?      �?433333�?�t�bj#  j�  j5  j�  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�C  j�7  �0.6�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�C  j�7  j�D  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubj8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C�������?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j3?  j[+  j4?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�K aj7  j�D  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jO?  j[+  jP?  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                       �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  ]�Kaj7  j�D  ��j	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jk?  j[+  jl?  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  j�D  ��j	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  j�D  j�7  �0.8�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj   hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  j�D  j�7  j-E  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubejG>  ]�j8  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        js+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jWE  j.8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  K j#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �       �       �              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�K aj7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jsE  jT8  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j18  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�Kaj7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�E  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K Kej7  ]�(K K ej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj-  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj4  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�8  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@333333ubaubj�7  G@      �_bounds�Nh��outward�G        ��j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C         ����p�        �J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ub�_patch_type��line��_patch_transform�j�  )��}�(h�}�h�Kh�hRh�Nububj�8  j/7  )��}�(h@�hANhBh�hChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  j;7  jK+  �jL+  j<7  jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jA7  jh+  jm+  jB7  j�8  jC7  jG7  j�7  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?����p�      �?�J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububj�7  j/7  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  j;7  jK+  �jL+  j<7  jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jA7  jh+  jm+  jB7  j�7  jC7  jD7  �XAxis���)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�	  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jR7  �jS7  �jT7  jV7  )��}�(j%+  j[7  )��}�(j^7  h7j_7  �j`7  Nja7  Kjb7  hhK ��h��R�(KK��h!�C(      �?       @      @      @      $@�t�bji7  hhK ��h��R�(KK
��h!�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�bjp7  �jC7  j F  ubj�7  j�>  )��}�(j�>  Kj�>  K j�>  �j�7  �j�>  �j�>  K j�>  �%1.0f�j�>  �j�>  j�>  j�>  �jC7  j F  j�7  hhK ��h��R�(KK��h!�C              9@      I@�t�bubj�7  �j�7  �ubj|7  jV7  )��}�(j%+  j�7  )��}�jC7  j F  sbj�7  j�7  )��}�(jC7  j F  j�7  hhK ��h��R�(KK ��h!�j�6  t�bubj�7  �j�7  �ubhchZ)��}�(h]]�j�7  ah`hbhc}�j�7  }�K j+  h�h�j�7  ��R���R�(j5F  h~��}�j�7  j�7  )��sNt�bssheKhfNhg��(K �ubj�7  �j�7  j�7  )��}�(h@�hANhBNhChGhIjS	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  h0h!C      8@���R�j�7  �Distribution�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@&      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  �top�j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�7  j�7  )��}�(h@�hANhBNhChGhIj_	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  h0h!C9��8�c9@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�7  G@      j
7  Kj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  Nj�7  Nj�7  �j�7  j�7  j�7  j�7  j�7  G?�      j 8  j8  )��j8  ]�(jD7  �XTick���)��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�	  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C        ���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�F  �_set_tickdown���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jrF  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C        �t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C                �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�F  �_set_tickup���R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jrF  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�F  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  jrF  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jrF  j�  K j�7  �0�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jrF  j�  Kj�7  jG  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNjC
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      9@���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j3G  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j$G  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      9@�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      9@        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      9@        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jiG  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j$G  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�G  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j$G  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j$G  j�  K j�7  �25�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j$G  j�  Kj�7  j�G  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      I@���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  jF  j[+  j�F  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�G  ��j7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�F  j[+  j�F  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�G  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�F  j[+  j�F  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j�G  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�G  j�  K j�7  �50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�G  j�  Kj�7  jQH  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubejG>  ]�jdF  )��}�(h@�hANhBh�hChGhINhJ�hK�hL�hMNhNj�
  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        js+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j{H  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�K aj7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�H  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�K aj7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj   hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�H  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K K ej7  ]�(K Kej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  Kj�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@333333uba�_tick_position�j�7  ubj�7  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C                 33333�F@        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�NububjNF  j/7  )��}�(h@�hANhBh�hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  j;7  jK+  �jL+  j<7  jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jA7  jh+  jm+  jB7  jNF  jC7  j F  j�7  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C               �?33333�F@      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububub�xaxis�j F  �yaxis�jG7  jV+  �white��_frameon���
_axisbelow���_rasterization_zorder�N�ignore_existing_data_limits��hchZ)��}�(h]]�(�xlim_changed��ylim_changed��zlim_changed�eh`hbhc}�heK hfNhg��ub�_xmargin�G?��������_ymargin�G?��������_tight�N�_use_sticky_edges���
_get_lines��matplotlib.axes._base��_process_plot_var_args���)��}�(�command��plot��_idx�K �_cycler_items�]�(}��color�G?�G?ܜ�����G?�TTTTTT��s}�j/I  G?�������G?�xxxxxxG?������އ�s}�j/I  G?�YYYYYYG?�G?���s}�j/I  G?䴴����G?�G?���s}�j/I  G?�������G?�������G?���s}�j/I  G?�G?�YYYYYYG?�[[[[[[��se�
_prop_keys���(j/I  �ub�_get_patches_for_fill�j&I  )��}�(j)I  �fill�j+I  K j,I  ]�(}�j/I  j0I  s}�j/I  j2I  s}�j/I  j4I  s}�j/I  j6I  s}�j/I  j8I  s}�j/I  j:I  sej;I  ��(j/I  �ub�_gridOn���_mouseover_set�hX�_OrderedSet���)��}��_od��collections��OrderedDict���)R�sb�
child_axes�]��_current_image�N�_projection_init�N�legend_�N�
containers�]�(�matplotlib.container��BarContainer���(j7+  j+  j�+  j�+  j�+  j�+  j,  j-,  jJ,  jg,  j�,  j�,  j�,  j�,  j�,  j-  j2-  jO-  jl-  j�-  j�-  j�-  j�-  j�-  j.  j7.  jT.  jq.  j�.  j�.  j�.  j�.  j/  j/  j</  jY/  jv/  j�/  j�/  j�/  j�/  j0  j$0  jA0  j^0  j{0  j�0  j�0  j�0  j�0  t�����}�(�patches�]�(j7+  j+  j�+  j�+  j�+  j�+  j,  j-,  jJ,  jg,  j�,  j�,  j�,  j�,  j�,  j-  j2-  jO-  jl-  j�-  j�-  j�-  j�-  j�-  j.  j7.  jT.  jq.  j�.  j�.  j�.  j�.  j/  j/  j</  jY/  jv/  j�/  j�/  j�/  j�/  j0  j$0  jA0  j^0  j{0  j�0  j�0  j�0  j�0  e�errorbar�N�
datavalues�hhK ��h��R�(KK2��h!�B�         @              �?              �?       @      @      @      @               @      @      @      *@      &@       @      &@      3@      4@      >@      :@      ?@      E@     �E@      >@      <@      4@      6@      =@      5@      2@      1@      ,@      (@      *@              &@      �?      @      �?       @      �?       @      �?                      �?              �?      �?�t�b�orientation��
horizontal�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�jZI  �remove���R�hQ�_container0��stale��ubj]I  (j1  j/1  jL1  ji1  j�1  j�1  j�1  j�1  j�1  j2  j42  jQ2  jn2  j�2  j�2  j�2  j�2  j�2  j3  j93  jV3  js3  j�3  j�3  j�3  j�3  j4  j!4  j>4  j[4  jx4  j�4  j�4  j�4  j�4  j	5  j&5  jC5  j`5  j}5  j�5  j�5  j�5  j�5  j6  j+6  jH6  je6  j�6  j�6  t�����}�(jbI  ]�(j1  j/1  jL1  ji1  j�1  j�1  j�1  j�1  j�1  j2  j42  jQ2  jn2  j�2  j�2  j�2  j�2  j�2  j3  j93  jV3  js3  j�3  j�3  j�3  j�3  j4  j!4  j>4  j[4  jx4  j�4  j�4  j�4  j�4  j	5  j&5  jC5  j`5  j}5  j�5  j�5  j�5  j�5  j6  j+6  jH6  je6  j�6  j�6  ejdI  NjeI  hhK ��h��R�(KK2��h!�B�        �?                      �?              �?      �?              �?      �?       @      �?      @      @              @       @      @      @      @      @      @      @       @      @      @      $@       @      @       @       @      @      @      �?      @      @      @      @      �?      �?              �?              �?      �?                              �?      �?�t�bjlI  jmI  hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�jZI  �remove���R�hQ�_container1�jwI  �ube�_autotitlepos���title�j�7  )��}�(h@�hANhBh�hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  �normal�j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ub�_left_title�j�7  )��}�(h@�hANhBh�hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G        j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�I  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ub�_right_title�j�7  )��}�(h@�hANhBh�hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�I  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ub�titleOffsetTrans�j�  �patch�j6+  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  jN+  jK+  �jL+  j7  jM+  jN+  jO+  jI  jV+  (G?�      G?�      G?�      G?�      t�jX+  G        jY+  K N��j[+  K N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  G        jo+  G        js+  G?�      jw+  G?�      j{+  G        j|+  j}+  j~+  G?�      ub�axison���	fmt_xdata�N�	fmt_ydata�N�	_navigate���_navigate_mode�N�_shared_axes�}�h�]�(h�h>es�_twinned_axes�Nube�artists�]��lines�]�jbI  ]��texts�]��images�]��legends�]��subfigs�]��suppressComposite�N�_layout_engine�N�_canvas_callbacks�hZ)��}�(h]]�(�resize_event��
draw_event��key_press_event��key_release_event��button_press_event��button_release_event��scroll_event��motion_notify_event��
pick_event��figure_enter_event��figure_leave_event��axes_enter_event��axes_leave_event��close_event�eh`hbhc}�(j�I  }�K �matplotlib.backend_bases��_key_handler���sj�I  }�Kj�I  sj�I  }�(Kj�I  �_mouse_handler���Kh�hG�pick���R�uj�I  }�Kj�I  sj�I  }�(Kj�I  Kh�hGj�I  ��R�uj�I  }�Kj�I  suheKhfNhg��(K KKKKKKK�ub�_mouse_key_ids�]�(K KKKKKKe�_button_pick_id�K�_scroll_pick_id�K�bbox_inches�j�  �dpi_scale_trans�hό_dpi�G@Y      j�*  hҌfigbbox�hҌtransFigure�hՌtransSubfigure�h�j�I  j6+  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  (G?�      G?�      G?�      G?�      t�jK+  �jL+  j�I  jM+  jJ  jO+  j�I  jV+  jJ  jX+  G        jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  K jo+  K js+  Kjw+  Kj{+  G        j|+  j}+  j~+  G?�      ub�_original_dpi�G@Y      �subplotpars�hD�SubplotParams���)��}�(j-7  G?�      j�7  G?�(�\)j�8  G?�������jNF  G?�(�\)�wspace�G?ə������hspace�G?ə�����ub�_axstack�hD�
_AxesStack���)��}�(hB}�(h>Kh�Ku�_counter�Kub�_axobservers�hZ)��}�(h]Nh`hbhc}��_axes_change_event�}�sheKhfNhg��ub�number�K�__mpl_version__��3.8.0�ubhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�hGh���R�hjNhkNhlNhmNhnhohphs]�]�����hx�h�j�  j�*  h�)��}�(h�}�h�K h�hRj�  hhK ��h��R�(KKK��h!�C       �?(\���(�?�������?)\���(�?�t�bj�  hhK ��h��R�(KK��h!�C      �      ��t�bj�  �j�  hhK ��h��R�(KKK��h!�C                       �?      �?�t�bubj�*  h7j�*  j�*  j�*  j�*  j�*  }�(h~�h��uj�*  Nj�*  Nj�*  h�j�*  h�)��}�(h�}�h�Kh�hRj�  hhK ��h��R�(KKK��h!�C �?IoN�?���`C!⿡�Wۦ@ڜ��H��?�t�bj�  hhK ��h��R�(KK��h!�C�?IoN�? �iK?�t�bj�  �j�  hhK ��h��R�(KKK��h!�C       �      �      ��      ���t�bubj�*  j�  j�*  jl  j�*  h�j�*  jt  j�*  h�j�*  h�j�*  j�  j�*  �matplotlib.gridspec��SubplotSpec���)��}�(�	_gridspec�jkJ  �GridSpec���)��}�(j-7  Nj�7  Nj�8  NjNF  Nj"J  Nj#J  NhChG�_nrows�K�_ncols�K�_row_height_ratios�]�Ka�_col_width_ratios�]�Kaub�num1�K �_num2�K ubj +  Nj+  j+  h�j+  j&+  ��R���R�(j~J  (K K KKt�}�}�j.+  h�j+  j.+  ��R�st�bj2+  ]�(�matplotlib.collections��PathCollection���)��}�(h@�hANhBh>hChGhIj�  )��}�(h�}�h�Kh�hRh�NubhJ�hK�hL�hMG?�      hNj�  hONhP�hQ�Train $R^2 = 0.885$�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j�J  �remove���R�hjNhkNhlNhmNhnNhphs]�]�����hx��_A�N�_norm��matplotlib.colors��	Normalize���)��}�(�_vmin�N�_vmax�N�_clip��j 8  NhchZ)��}�(h]]��changed�ah`hbhc}�j�J  }�sheKhfNhg��ubub�_id_norm�K �cmap�j�J  �LinearSegmentedColormap���)��}�(�
monochrome��h8�Greys��N�M �	_rgba_bad�jN+  �_rgba_under�N�
_rgba_over�N�_i_under�M �_i_over�M�_i_bad�M�_isinit���colorbar_extend���_segmentdata�}�(�red�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�green�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�blue�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?�?�?      �?;;;;;;�?;;;;;;�?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?�������?�������?      �?                �t�b�alpha�hhK ��h��R�(KK	K��h!�C�              �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?�t�bu�_gamma�G?�      ub�colorbar�NhchZ)��}�(h]]�j�J  ah`hbhc}�heK hfNhg��ub�_us_linestyles�]�K N��aj�6  ]�h0h!C        ���R�N��a�_us_lw�hhK ��h��R�(KK��h!�C333333�?�t�b�_linewidths�j�J  j�6  N�_face_is_mapped���_edge_is_mapped���_mapped_colors�NjI+  jJ+  jO+  hhK ��h��R�(KKK��h!�C �?�������?TTTTTT�?      �?�t�b�_facecolors�hhK ��h��R�(KKK��h!�C �?�������?TTTTTT�?      �?�t�bjL+  �face��_edgecolors��face��_antialiaseds�hhK ��h��R�(KK��h�b1�����R�(K�|�NNNJ����J����K t�b�C�t�bj
7  G@      �_urls�]�Naj`+  Nj�7  Kja+  Njh+  N�_offsets��numpy.ma.core��_mareconstruct���(jK  �MaskedArray���hK ���b�t�R�(KMK��h!�B�!  ޯuŢ��?��m��������?�$�޻ۿ6Ah"���?�	B��?K�C.���?��'�3-���i�`��?�@'���?� �����? �H�?��AU�@��d/�����Az4@@e�Շb�����w��? l�Cy;U?�Hc�pw�? �c�ޭ�W�$K�!�?�ڵM�罿��_��? ����n?���@�l9�*�?sgn����?�;sSu�?IJɧrB�?X\X��<�?8���Y�@@Aߓ���?�� ,�@`j�Lg���h�Ҧ�?��]�?��>�1�?�#Z�?��.�zB ��?��=4��?<����@@l�a�����S��v@��[+����L3�? }�f���?n��`�i�?P�y$���6�>�$�?��+��?�0�@�r�����?,�+��� @8P:ӿ�e^��`�?�ړ�p�Qh��@@��G�_�?~A��@P�U��� %�ߩ@ �f�/F�?�w���?P~��vmȿ��|����?�ǆ�Nǖ?rB!���?�����ĵ��Xd}0�?��E�ð?�n�Lq�?H��#�?I��uY�?th��3\ٿ�N��9��?h��p0vȿ9�J���?`��u\Ơ?틞�d��?@k�0&�?�P��*�? BM<ª�?�bf�?p�!6Aa�?��n=�@ ���¥?�y�ث�@ F_N�v�s9��Z��? 8?�{���ˮt���?x�D-f пf�,]oA�? ��{��r��%|@ �~����K���\+�?�q�Y���?"���@@��ɫ��p�S��?����:������</�? �[�L������Dv��? ]V&�+�?�hL���?(�:��ܿ�Iȷ;�?����A"οhp �,�? ��2�1��|aA�\��?�:A	n���)ᔒ'�@���'���hze��?����A���g.��?0��[�ο\�Q"җ�?`����?~%O�@�W�$��?3�W���?��'��m�?�W飩@ � �-��?�O֔$@��#Z4,�?/h�5��?�&Z�?c=m_z�? ����s?=��#"�?@
�������0^�? mGKࢪ�1/�+��?Ps��뵿�՜�E@ ��0����B4i���@�`ll�?XӮ}JS�?@�邜�?�ܻ�'f@ iH̑�?��T�f�?H�8�B5�?�,�!��?�e�&1�?w�:��?'�:��?��#�{��?��G��$�?�5�ܜ�?xH����?屄�֔@`	c]�g�?G{	���?�@��u��?�����a�?����E׿U3V@&��?1at���d>��?�K%�r��p���w�?`ؒ�t��E�x�iN�?���@�?xY�9�?��ڈ��?�-Nڐ��?���ɿ?�[i3us�?\]'���ֿ��NȢ�?�t���?�guB��? *J���?�/M��.@��r���?������@ Z�
���?����
 @ ����
�?Y�@@���6��mN�s$��?ڜ��H��?>S�ܺ��?�35ȭ��?|�w�h�?@xĎ�v��J�T����?�yo>Fҿh����?�{;��?���>
�?D��\�������@�Q��L�?B'�� �?�&q���?"(�R|H�?����?D+��H�?� Z�D�?2��Ta��?��c�@ӿ�x�&���? Y49_��?��'2'@ >�\x�~�޷�` @�_��-5�?$N��q�? ��nk@�?�=u���@ +]a�n���9l�?P,��o���$���?1�V�ɿ�7�>� @���}RǿS�(#I @ /R��P׿DU,F�a�? �D耤Q����".��?�p|�zؿ".Y���?�q���?�sR�?�?��؊����9�D�@ ��O$��?�ǇPy��?`�ӻ�]���8ҵ��?��q|����2����?�^!�{ټ?�7��a�?`#z��i�?ni�8#� @�-�g��?׉:��@ �xP��?��=�Rt�?���<N�ӿ�2����@��Г���G��h�@ ��5e̕�e�ޡ�d@�{�{z���A��~+�?���{�=ȿt�},t#�?`��^�οnH���,@ K�,0���'���:�?��m�RS��������?���1��¿��-;P��?�M��ݿ��\�&�?P�����?��/>�?���O�οv��1
@ w@��?��%�E�? ���r?�X%� ��? ��D�?�A9�W�?H�I���?#��I�?趓�%ϿMd��p�?�Έ���?��c��@�`�&Z����i��@ I�We%��u3xÄ�@��_�͕��@�����@�a��9��?�u��x@��83wȿ��},K@ ��},K�?Zl�J�E@ P��뤿�^07J�?��s��?�u�tڄ�?���b�ڿC>�Tz��?���x�jڿ.`s�+@(��e!:п[�)L���?��.w��?.4 ��B@@z�߈������2p��?@���?�?���pm@�s�Y����qX��?���ú�? 1��'&�?�������?�3��?�Kl\�����i¿?�?Ppe}b�?&4���V�? n.����?8H���@ }�AT�?$g�Ku�? ��q�����c�@0��VͿz�67�?�O��?�T
�?(��z�Կ����� @�}���?�W<�d�?�U4z���?(|�W[��?`�Mܾ~̿��b,�@_�-ƒ�?i �U���?��(P�������Y�?��+:�0�?[D�I�?@H�[d���Q��&�?���U4пH�3�; @��`�ſs�{u�@ [6����?�6~vnT�?@k�g�F�?����@�,�)'�?�1�?x��p���?a�. � @ �c-���ȯ�F��?����?��<�+d�?��L����0�@���MnӤ������B�?���B�>�?�]�r�@�<��'�?Ă�I���?���x��?Q�飩��?ŝ>�z�?���_��@@�Kq�?]w�y @ �ݼ\���l�:�j�?`��C}D�?������?X��U%O�?��t�U�?�h蠒�?J=�S���?����?k����r @�J=�j¿����ʯ @�4}��9��R�L��? ��Ks���O�^:���?�>�?]e�?$=x��o�?�`��e6��Q'���� @ In�"��l�A\�? ��F��?�9@�!b������
��?8;��^�?7��kQ�? ٬��ݥ�4��u@���F�ޑ�8�뉐�?���j������@��R �S����b�]�@`y�eU%�?B�L�8e�? @��2����-��?�Y�TP����o+@�E,h��Ŀ�簮�?�E۷G��?���}b�@  ���\�4�K���?�?���G��xWxY���?�����8����f�P�?���7��?����\@PL���Z�?�&IzD�@ Pٶ����h�͙���?��[Y&_��W/>K��?�#_s�C�?0_���@��_���?	��0��?Ȋ"�(�?�d�8]@�����?�x�3��?p�%�ּ�?0��!���?b�"И�{ U�v��?`�(��ݧ��������?���T�f��WRr+��?���`C!⿤��]�?�X�U��wT�a��? ��<�~�s�o9'��? :�1���?�I��?�ǁu���q\e���?�>!��i��!� �D�?	�%�?n(܍q@@�zD�Q���!A���?0��˿˾�&+ @��8�ƿ6F���? ���ݔ�ݾe�0~�?O�j�ٿ�n�Ѧ�?xu�'�6�? ��^��?�,�����ˁz�?��T�A�?هt�K��?�RbT�?:���S�?0�Rgſo�Fq�? ~V1�e?~*=���@���ɘ�?h��b�O@ Z����?v�)��@`(�^xs�?��j���?`��I�A�?�2�zLH�?���$ĿrG�%���?@���'��4��i��? gJU���?�`�\-�?�J�Y�Կ��GX�-�?��?��l�?�a}�ݝ�? 0��������o!���?��qoJ�?����F @ =��1��?kP�PS�?��+�+&п�
�#�q@ r�YH����oH�@����@�?���!�$ @��:b�����mӐ�@�S�R�?�Rx׷�?`s��?/�	n@���G?��	�� @@8��#��?���e���?�0p����3�3!��?�������L(E���?������J���e@�v|(@B���}��ޔ�?��^AQyҿ"��/��?@t�i#E��p>=���@ ��c���?ȟM�"��?@�l���?^�b���? Q��N����#�?��??R����?���~��?��%b>�?QDZ@�c���?l�)^}l�?cu{ÿwm�d��?�� ������v[��?Щ�{]����.����?�o��X��?@�Y闧�? 0+��?l
8����?|��uO��?$�w��=�?� �;Y�����=�'�?��5iR��ϴui�� @p�ʿ"��_l @����%��c�:(�?D���,Կ���~@�5��rC˿����G4�?��e>����"^��b�?����?>��K��?���]��?}}�8ą�?���kA��?����?���ڳ��?�j�?��?@�|:�h��O�����?L1�Q&�?l�d�!�? :GFtп�n%m��?�tC(i��?��[���? �k��aT���g,$x�?@i��a��z��Tf��?��Ke�?��8��?��O�>ӿ�q�q"�? �5iDi�?<W�H1@�����Qÿk�5�
��?��#���?,��RG�@��m.u�?,��7KT@����D�?�)����?�Tߗ˚���p<@�? J���Ϝ?�Q	��?���!�A�?(=�����?@�D�?�ǳ��^�? �y��]��>4Y�#�?b7�S��?�k��@ �k�ă?��/�� �? ���<��*-P�e�?H�0jƿ*Qz���? kW�¶v��[w�Ek@��*��>�(���?����{���ǁ�D@@�o����2���?`g�<c(��:XJK���?`q��8�ÿ��:���?H=�ǂ�Ŀ��B=��? T;��v�@%|b���?h�V��?R��B�@��ǧ��?eM0%a�?`�\�Yۣ�$~F�׿@�C-{�֬�MB�rT��?0��Ŀ$���@ yF+:��[lJ�U�@`A¶���Xb�@`t���е���kRp@P�s|.̿*3����?��03���?�l���?`���힤?!y�m�@H^����п���I���? ��nظ���!;@���q.�?�S���?��}/�?R�N�;��?G�uO������w�?��Vt��x��J�W@���h����=�J�@@i����hf��>O�?���2 '�?^*�[�?x��o=H�?] {����?��qMg�?���w�4@�v�H��?1��z!}�?�!����?��|",� @ w�>��Ϳ��2�@�2�������!�=�?�I�AZ���A�A��@�Y�N�뮿����@��? L/Խ?%�&�@�X��(�?V	D�TF@ #�V!�?r��U�?P
��(��?+��O��?��f�?��?)4��g�? {�t�Q�?Hv6][��?���_}�����v��i�? �iK?��F���?���7R�?�Q����@�����?�n���@ �x0��?LRt�,��?�9�o����cx۳��?��Y��/�����s���? k�:���?�������?��7t=$�?�/����?�K�C��?�=$ny�@@$�i�ƿxMiA���?�kJe�?j(,=��?��p`�ò��4M����?��i��E�?z߅��?�Eu޽�(V��s��?`�f��-Ϳ���8ʦ�?@�HK��������\�?@
gj�ɪ���,�Z�?T����.п��vi��?`+b�Ʀ?���ٔ @h�)��Կo>n �@�jRjC@�?����b@ {�w�a��1Y�ۂ��? c�w��?DU��V�?x������?K.:�v�@��3nw�?(:N���?�.>��˿�C��)�?�E� ޴�?��_���?�AZ�| �?h�Y�,�@�&��.��?������?�?F08���H�D�?�%^#ڽ?CANsv��?0�4g׾?�"v����?@(b����?W��X�?�E/��S�?vʇ���@ AR�E�?x���3@��-ÿ��U��R @ O=�nĿh��E�?@k��p,�?U׶�?�5k��?���R��@����ִ���Ǒ����?����ڿ%�S���@����?z���P@ ���E����x��?�T~T�>ڿh���Hp�?8J�O�?���D�?�ê��&�?n��(�? ��bJaf�*��`�@@<��_��?�Y��^�?t����?���>D�?p���?��� ��?`�a�?<��(���?P-�i#ǿ��,�ݶ�?@�e<v�?DX�;�2@ �wm�{����ҏ@ Z��K���{���@�Z{8�S�?~>���@ ��kQm�����L�}�?Ȝ5�ſ���_��?�g&l���a}C��?�xWA�ț�-d��|�?����Ŀ��0�ێ�?@����?���$\�?�S���q��T�%��?�k8-v=���u}�e�?�[�p���?��@���Y���?qY@�q�? ��De?��b��@�|�y@JM�4@�?`����ѧ���tߴF�?HiXY�ſ$֠㩽�?�C��Sb��GP�uA��?�^��Ͳ?)8gL��?Rp��$�?�U�)�@��-���?��i�@��/�׿������? �I�cS��T,6t�@��AH�/���h�LHA@ �j�2*|?K��Q���? �e�Dx�ko_�C@�����
�?>��	dg�?���Jy^ο���I@ ���|M�?0��q@ ����=�����c��?��3�狿P�SY$R�? wBt�����d�?�=�a��?�`:��i�?P�,6�Ŀ*���-�?P�Twdn�? k����?�@F-:	̿�n����@ ������?��")���?��I��?��,��@@������?��(2��?`�	ſ~����?���ڞ��?�󚩭�@�^#��Q�?�"�,O�?p,2���?�P�(�@�E����?�~�NL�?�A,p%v���# �b�@�Ko�"?�?v��)�P�?�]�m�+�?`b#��@ &6R���?C|ޢC�? �I�op?���6�p�?�S\́�?�aP3�?�1��Ԍ��A�����?�=����¿ze� ��?�s��Hנ?���|H�?�$}͉��?��#����?�&-�[���'�o�? 
��a��ҕ,���?�S,tܦ?��^z7@�jy���¿g�L�־�?�l��H	ʿ;a1�[�?=���?���"1�?p�
$^�?Vz@��6�? �G����Ew��/�?��6bMԿ\���@ ��i�m?Ch��c��?`��q��?CW8�7d�?���'�wοNɹ-��?t8%�x�?j�p���?���\_K��B��j�@��:0��?���2���?��k�����p�O�E�?�	����ӿڄ�n�@�4J�[��?l�І @8c�xٿZjN��)�?�F&/�Lȿ�+C��?����ѿ7|����?��S�<��?��
���?���Jc��$�wP�&�?�P��?�����M@�:��5��?�4M@ G��^��%��?� �M
t��N���	@�p�ܽM�?3�e�@ �J��C�-���? ��l��r��Aɢ�@����?Zi�@���?`j��˦���2��?���9�í�������?@�Z�	w��6-:��?���T �?��,K�@@foeY��?���{���?��T��ÿ �Y�@ �Qg�_ƿ`�2���?0-�CQ�����Zs�?;�<���?1O�ν��?��^�ve�?�%pz�?���2����K��?@z>���DM6���?@$�2����Բ4��?�������?��ƅ��?�����5�����Mr�@��U�x��nޭ0���?p�n��^�?t:E4z�?�O��Ȱӿ̦�53w�?@c����Ϳ�����@ � !�����#f$��@��C�Щ��N�[t��?�%w���̿����@��A���п���G�? �q>P���^|$���? ~�ol��?;.I\m�?@�_�H��?+'�v� @`�$���?|z3V[
�? ,dN%���V!��@ �K�?�iJaP�?Ps��-��"-;�U@ q2��?"u7�k�?�(�E�Q��T�Zz�	@ ����s?�j��/ @�C�iaؿj��w�?��?��辿
��=I�?�Ba�@O�?�)��H$�?@3��i����s�2� @`���l��Uh�\�(�?`��aT꪿���%�? Rc�o&��4B���?��/"���B8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �Nt�b�_offset_transform�h�_paths�j&  )��}�(j)  hhK ��h��R�(KKK��h!�B�                �rSl��?      ࿉��e��?���֠ܿ�;f���?�;f��ֿ���֠�?���e�п      �?rSl���      �?              �?rSl��?���֠�?���e��?�;f���?�;f���?���e��?���֠�?rSl��?      �?              �?rSl���      �?���e�п���֠�?�;f��ֿ�;f���?���֠ܿ���e��?      �rSl��?      �              �rSl������֠ܿ���e�п�;f��ֿ�;f��ֿ���e�п���֠ܿrSl���      �              �              ࿔t�bj0  hhK ��h��R�(KK��h�u1�����R�(KjK  NNNJ����J����K t�b�CO�t�bj1  Kj2  G?�q�q��j3  �j4  �ub���_sizes�hhK ��h��R�(KK��h!�C     �H@�t�b�_transforms�hhK ��h��R�(KKKK��h!�CH�q�q#@                        �q�q#@                              �?�t�bubj�J  )��}�(h@�hANhBh>hChGhIj�  )��}�(h�}�h�Kh�hRh�NubhJ�hK�hL�hMG?�      hNj   hONhP�hQ�Test $R^2 = 0.895$�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j�J  �remove���R�hjNhkNhlNhmNhnNhphs]�]�����hx�j�J  Nj�J  j�J  )��}�(j�J  Nj�J  Nj�J  �j 8  NhchZ)��}�(h]]�j�J  ah`hbhc}�j�J  }�sheKhfNhg��ububj�J  K j�J  j�J  )��}�(j�J  �h8j�J  j�J  M j�J  jN+  j�J  Nj�J  Nj�J  M j�J  Mj�J  Mj�J  �j�J  �j�J  j�J  j�J  G?�      ubj�J  NhchZ)��}�(h]]�j�J  ah`hbhc}�heK hfNhg��ubj�J  ]�K N��aj�6  ]�h0h!C        ���R�N��aj�J  hhK ��h��R�(KK��h!�C333333�?�t�bj�J  jpK  j�6  Nj�J  �j�J  �j�J  NjI+  jJ+  jO+  hhK ��h��R�(KKK��h!�C �������?xxxxxx�?�������?      �?�t�bj�J  hhK ��h��R�(KKK��h!�C �������?xxxxxx�?�������?      �?�t�bjL+  �face�jK  jK  jK  hhK ��h��R�(KK��jK  �jK  t�bj
7  G@      jK  ]�Naj`+  Nj�7  Kja+  Njh+  NjK  jK  (jK  hjK  jK  t�R�(KK�K��h!�B�  ���X6
�?���G��L�f�w�@ �m��?Ay���)@���I��?y����? J��z��?���2�@�Gх������~���?h��p� Ͽ\���h�@�u껌�?�?IoN�?��M:�/ڿ�����?@I�}?[ܚ���?�>I=��? ��-���? `|o���?35h�}�? �_�<V��m�a���? �A�e�W?�&�e-1�?@)�MSڙ���Wۦ@�&�G�:�?�,��%��?��qZ�/�?�yX?@ ����t¿`s�,FS�?`0Ϛ2�����+@ �WA+��L䣓B~�?@F,�Ò?8G��5@��~��/¿�0�֌@�?��I�f�?��	�#��?h[���F����0��?���C9t�?���) @ x���?��=���? �4Jn��.	
H��?pIP@��?O�j ��?��0�i��?>Hy��? |kȂ﾿������?����j�ѿ�
��9��?�޲�c�ÿ�~�-��?��`�#�?�}E���?�r�)��?��c�c� @kz�}տ��3sA��?������̿*\���k�?�m:0�̿�K6�v@ 9������:�Ӷ��? u`Jԑ?���t�@��E!��ſ�$49� �?�$�"]��а~�.R@ �7�"�?�׊��v�? }�8Jo�?��W��k�?��`��L�?.u_d��?Pn+��?�_�
�?�2��U��?��o���?P����?���l��@���Φ��?U�3Ĥ�@ "YF48��@�c��E�?�?>ҵӿT�3���@��Ԭ���?�J�F�@��}�]��$��Rsr�? )|����?vIP�7�? b<=,��?�����%@���ns�? M��&�? hj��4�?!�;�NJ�?���$Gǿ���YB@��Q�l���0;��N�?(Sk ���?n�>�?�a��?	ٸ�?�?X�һ��Ͽ�c�
 @\���ȿZ^Y3�@@6u��?��m�x�+�?���N�����"�,@@�fi��?E8ڡ� @�=,��ؿ�p�X@`*��ĪͿ��Z���? �X�v��K��e�i@ AP�e�?��`v҇�?`�Ll�ÿ�ޣ��? ���Y+�?�i��@ x�*p�?�Ő��@P�&J�ƿ9��@@�#�Q�?�!Z�[@ ]�� ���YQ�F�?���ɾ�W���N�?�{25v���������?��5�����)�����?Г���״���Ҧ|:�?�P�������~z@HM����? ���@��B{�8�?[d�I��?X��ÿ�������?�Ҍ:��п�J9+d�?�֘z��\'���@ ��nS��T�Z��? ���<z�?&0�+�-@ 8���?ta}��@�ot�i˦�zX�t�?�:��?S��,d%�? �-�k�7���/@�S�%�˲?2�㮅�?(k���?F�璣�@��唟��?����)��?�<�N��?`>�j��? 4���A��v��ψ@����f�?k��ȸ@ �1k�.�?�����5�?�44�����Z����? w��Œ�? �JEf @ i��̂��N%�<��?�t*��I�?��&�ʈ�?��S�?D��e'�?�~-J��M�_�$@ ��K�|�1.R����?P�Ca���R���? �N)Ȃ�?�=�M�?�w�nb�?vc�X]@�����?��{��?���U�?«#Ĕ��?P�mu��?�>��1��?0G��@���T�%@�y�%�ĿY�B��?H/Q�|(�?�D��@ d��-�?������@ V��0��?z��ϫ�@����YпLJ�����?��l��?0����s@���X���?� �:� @`Y��Rǿ�?����?��P6��?�կ��@��c� ���x��L�&�?@b���?���
��? a�I���?���	_�?`~��ɑ�?ƿ��I�@ �I�l�?q-EP�? \�~�1��@{M�	�? e���ʵ���Z,��?�Ōa�ѿ*yz`r�?(�R�J߿�H��I��?`Q=,��� �S�@�][$��?�Q��S@� �o�������@��j[2׿�UN����?@��-��?Gi�p�?��ѯV?����-^���?��%����B                                                                                                                                                                                                                                                                                  �Nt�bj#K  h�j$K  j&  )��}�(j)  hhK ��h��R�(KKK��h!�B�                �rSl��?      ࿉��e��?���֠ܿ�;f���?�;f��ֿ���֠�?���e�п      �?rSl���      �?              �?rSl��?���֠�?���e��?�;f���?�;f���?���e��?���֠�?rSl��?      �?              �?rSl���      �?���e�п���֠�?�;f��ֿ�;f���?���֠ܿ���e��?      �rSl��?      �              �rSl������֠ܿ���e�п�;f��ֿ�;f��ֿ���e�п���֠ܿrSl���      �              �              ࿔t�bj0  j/K  j1  Kj2  G?�q�q��j3  �j4  �ub��j8K  hhK ��h��R�(KK��h!�C     �H@�t�bj?K  hhK ��h��R�(KKKK��h!�CH�q�q#@                        �q�q#@                              �?�t�bubj�6  )��}�(h@�hANhBh>hChGhIj�  hJ�hK�hL�hMNhNj^  hONhP�hQ�_child2�hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�j�J  �remove���R�hjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j�6  j�6  j�6  )��}�(j�6  h�j�K  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  j�6  j#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j	7  �j
7  Kj7  K j7  ]�(K Kej7  ]�(K K ej�  hhK ��h��R�(KK��h!�C              �?�t�bj�  hhK ��h��R�(KK��h!�C                �t�bj7  hhK ��h��R�(KKK��h!�C                       �?        �t�bj#  j�  j5  j�  j#7  �j$7  Nubej%7  ]�j'7  j*7  )��}�(j-7  j/7  )��}�(h@�hANhBh>hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  j;7  jK+  �jL+  j<7  jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jA7  jh+  jm+  jB7  j-7  jC7  jq7  j�7  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C         ����p�        �J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububj�8  j/7  )��}�(h@�hANhBh>hChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  j;7  jK+  �jL+  j<7  jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jA7  jh+  jm+  jB7  j�8  jC7  jq7  j�7  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       �?����p�      �?�J�Qv��?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�Nububj�7  j/7  )��}�(h@�hANhBh>hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  j;7  jK+  �jL+  j<7  jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jA7  jh+  jm+  jB7  j�7  jC7  j�E  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jR7  �jS7  �jT7  jV7  )��}�(j%+  j[7  )��}�(j^7  h7j_7  �j`7  Nja7  Kjb7  hhK ��h��R�(KK��h!�C(      �?       @      @      @      $@�t�bji7  hhK ��h��R�(KK
��h!�CP�������?�������?      �?      �?      �?       @      @      @      $@      4@�t�bjp7  �jC7  jL  ubj�7  j�>  )��}�(j�>  Kj�>  K j�>  �j�7  �j�>  �j�>  K j�>  �%1.2f�j�>  �j�>  j�>  j�>  �jC7  jL  j�7  hhK ��h��R�(KK
��h!�CP      �?      �?      �?      �?      �?      �?       @      @      @      @�t�bubj�7  �j�7  �ubj|7  jV7  )��}�(j%+  j�7  )��}�jC7  jL  sbj�7  j�7  )��}�(jC7  jL  j�7  hhK ��h��R�(KK ��h!�j�6  t�bubj�7  �j�7  �ubhchZ)��}�(h]]�j�7  ah`hbhc}�j�7  }�K j+  h�h>j�7  ��R���R�(jCL  h~��}�j�7  j�7  )��sNt�bssheKhfNhg��(K �ubj�7  �j�7  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  h0h!C      8@���R�j�7  �Predicted Value�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@&      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�7  j�7  )��}�(h@�hANhBNhChGhIj�  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  Kj�  h0h!C9��8�c9@���R�j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�7  G@      j
7  Kj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  }�(j�7  �j�7  �j�7  �j�7  �j�7  �uj�7  Nj�7  Nj�7  �j�7  j�7  j�7  j�7  j�7  G?�      j 8  j8  )��j8  ]�(jdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNjR  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�L  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j}L  ��j7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�L  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j}L  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�L  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j}L  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j}L  j�  K j�7  �0.50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j}L  j�  Kj�7  j�L  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jM  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jM  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jPM  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jM  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�jlM  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  jM  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  j'  j5  j   j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jM  j�  K j�7  �0.75�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jM  j�  Kj�7  j�M  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�M  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�M  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j�M  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  j>  j5  j;  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�M  j�  K j�7  �1.00�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�M  j�  Kj�7  jJN  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R��a�      j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jgN  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jgN  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  jgN  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  jM  j5  jJ  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jgN  j�  K j�7  �1.25�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jgN  j�  Kj�7  jO  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jO  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jO  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  jO  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  j\  j5  jY  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jO  j�  K j�7  �1.50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jO  j�  Kj�7  j�O  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      �?���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�O  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      �?�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      �?        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      �?        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�O  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j�O  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C      �?      �?�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       �?              �?      �?�t�bj#  jk  j5  jh  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�O  j�  K j�7  �1.75�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�O  j�  Kj�7  jrP  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C       @���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�P  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C       @�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C       @        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C       @        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�P  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j�P  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C       @       @�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C        @               @      �?�t�bj#  jz  j5  jw  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�P  j�  K j�7  �2.00�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�P  j�  Kj�7  j*Q  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      @���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jGQ  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      @�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      @        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      @        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  jGQ  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  jGQ  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C      @      @�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       @              @      �?�t�bj#  j�  j5  j�  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jGQ  j�  K j�7  �2.25�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  jGQ  j�  Kj�7  j�Q  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      @���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�Q  ��j7  ]�K aj	7  �j�  hhK ��h��R�(KK��h!�C      @�t�bj�  hhK ��h��R�(KK��h!�C        �t�bj7  hhK ��h��R�(KKK��h!�C      @        �t�bj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C      @        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�Q  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j�Q  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK��h!�C      @      @�t�bj�  hhK ��h��R�(KK��h!�C              �?�t�bj7  hhK ��h��R�(KKK��h!�C       @              @      �?�t�bj#  j�  j5  j�  j#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�Q  j�  K j�7  �2.50�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�Q  j�  Kj�7  j�R  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubjdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  h0h!C      @���R�j8  �j�7  G        js+  G?�      j8  G@      j8  j�6  K ��j8  G@ z�G�j8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�R  ��j7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�6  )��j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C        �               �      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j�7  G@ z�G�j
7  Kj7  K j7  j�R  ��j7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  j�L  j[+  j�L  j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�6  )��j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubhIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  j�R  ��j7  ]�(K Kej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�R  j�  K j�7  �2.75�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj	  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  j�R  j�  Kj�7  j<S  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@      ubejG>  ]�jdF  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNjf  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j8  K j8  �j�7  G        js+  G?�      j8  G@333333j8  j�6  K ��j8  Kj8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�jfS  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                       �      �       �                      �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�K aj7  ]�K aj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  NubjD8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j+8  j�6  �j�6  j�7  j�6  j�6  )��}�(j�6  h�j�S  j�F  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  Kj#  j�F  hIh�)��}�(h�}�h�Kh�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubj�6  Nj�6  Nj�6  G?�      jh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G        j_+  �j7  j�7  j7  G?�      j7  j7  j7  j7  j
7  Kj7  K j7  ]�K aj7  ]�Kaj	7  �j�  Nj�  Nj7  Nj#  Nj5  Nj#7  �j$7  Nubjb8  j�6  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMG?�      hNj�  hONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�6  jg+  j�6  j�6  j�6  j�6  j�6  j�6  j�6  Nj�6  j�6  jX+  G?�      jY+  K N��j[+  G        N��j]+  j�6  j�6  �j�6  j<7  j�6  j�6  )��}�(j�6  h�j�S  j�6  ��R�j�6  Nj�6  Nj�6  Nj�6  j�6  j�6  hRj#  j�6  hIj�  )��}�(h�}�h�Kh�hRh�Nubj�6  Nj�6  Nj�6  Njh+  j�6  ja+  jg+  j�6  �ubj�6  Nj 7  Nj7  G@      j_+  �j7  j7  j7  G        j7  j7  j7  j7  j
7  Kj7  K j7  ]�(K K ej7  ]�(K Kej	7  �j�  hhK ��h��R�(KK ��h!�j�6  t�bj�  hhK ��h��R�(KK ��h!�j�6  t�bj7  hhK ��h��R�(KK K��h!�j�6  t�bj#  j&  )��}�(j)  hhK ��h��R�(KK K��h!�j�6  t�bj0  Nj1  K�j2  G?�q�q��j3  �j4  �ubj5  Nj#7  �j$7  Nubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  jNF  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�7  )��}�(h@�hANhBNhChGhIj  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  Kj�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�8  j�8  j�8  G@333333ubaj�H  j�7  ubj�7  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C �Ԓ.�p�?        �[8^@        �t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�NububjNF  j/7  )��}�(h@�hANhBh>hChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  j;7  jK+  �jL+  j<7  jM+  j;7  jO+  j7  jV+  jN+  jX+  G?�      jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jA7  jh+  jm+  jB7  jNF  jC7  jL  j�7  G@      j�E  Nh�j�E  j#  j&  )��}�(j)  hhK ��h��R�(KKK��h!�C �Ԓ.�p�?      �?�[8^@      �?�t�bj0  Nj1  Kj2  G?�q�q��j3  �j4  �ubj�E  j�E  j�E  j�  )��}�(h�}�h�Kh�hRh�NubububjI  jL  jI  jq7  jV+  jI  jI  �jI  �jI  NjI  �hchZ)��}�(h]]�(jI  jI  jI  eh`hbhc}�heK hfNhg��ubjI  G?�������j I  G?�������j!I  Nj"I  �j#I  j&I  )��}�(j)I  j*I  j+I  K j,I  ]�(}�j/I  j0I  s}�j/I  j2I  s}�j/I  j4I  s}�j/I  j6I  s}�j/I  j8I  s}�j/I  j:I  sej;I  ��(j/I  �ubj=I  j&I  )��}�(j)I  j@I  j+I  K j,I  ]�(}�j/I  j0I  s}�j/I  j2I  s}�j/I  j4I  s}�j/I  j6I  s}�j/I  j8I  s}�j/I  j:I  sej;I  ��(j/I  �ubjII  �jJI  jLI  )��}�jOI  jRI  )R�sbjTI  ]�jVI  NjWI  h=}���jXI  �matplotlib.legend��Legend���)��}�(h@�hANhBh>hChGhIj�  )��}�(h�}�h�Kh�hRh�NubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhih�h>�_remove_legend���R�hjNhkNhlNhmNhnhohphs]�]�����hx��prop�j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ub�	_fontsize�G@$      j�I  ]�(j�7  )��}�(h@�hANhBh>hChGhIh��CompositeAffine2D���)��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}�����Hj6T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?-؂-��{@                      �?�t�bubh�h�)��}�(h�}�����Hj6T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?-؂-��{@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  j�J  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�7  )��}�(h@�hANhBh>hChGhIj5T  )��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}���r�Hj^T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?"""""Rz@                      �?�t�bubh�h�)��}�(h�}���r�Hj^T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�hhK ��h��R�(KKK��h!�CH      �?        @�~&f|@              �?"""""Rz@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  jKK  j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@$      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ube�legend_handles�]�(j6+  )��}�(h@�hANhBh>hChGhIj5T  )��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}��М��Hj�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH��8��8�?                        ��8��8�?                              �?�t�bubh�h�)��}�(h�}��М��Hj�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        \����y@              �?-؂-��{@                      �?�t�bubh�hhK ��h��R�(KKK��h!�CH��8��8�?        \����y@        ��8��8�?-؂-��{@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQj�J  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  (G?�G?ܜ�����G?�TTTTTTKt�jK+  �jL+  jK  jM+  j�T  jO+  jK  jV+  j�T  jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  G�       jo+  G�       js+  G@4      jw+  G@      j{+  G        j|+  j}+  j~+  G?�      ubj6+  )��}�(h@�hANhBh>hChGhIj5T  )��}�(h�Kh�Kh�}�h�K h�hRh�Nh�h�)��}�(h�}���v�Hj�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH��8��8�?                        ��8��8�?                              �?�t�bubh�h�)��}�(h�}���v�Hj�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?        \����y@              �?"""""Rz@                      �?�t�bubh�hhK ��h��R�(KKK��h!�CH��8��8�?        \����y@        ��8��8�?"""""Rz@                      �?�t�bubhJ�hK�hL�hMNhNNhONhP�hQjKK  hSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  (G?�������G?�xxxxxxG?�������Kt�jK+  �jL+  �g�jM+  j�T  jO+  j�T  jV+  j�T  jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  G�       jo+  G�       js+  G@4      jw+  G@      j{+  G        j|+  j}+  j~+  G?�      ube�_legend_title_box��matplotlib.offsetbox��TextArea���)��}�(j�7  j�7  )��}�(h@�hANhBh>hChGhIj5T  )��}�(h�Kh�Kh�}�h�Kh�hRh�Nh�h�)��}�(h�}����Hj�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�h�)��}�(h�}����Hj�T  sh�K h�hRh�Nh�hhK ��h��R�(KKK��h!�CH      �?                              �?                              �?�t�bubh�NubhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  K j�  K j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubh@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�j�T  a�_offset�K K ���offset_transform�j�T  �_baseline_transform�j�T  �_multilinebaseline��ub�_custom_handler_map�N�	numpoints�K�markerscale�G?�      �scatterpoints�K�	borderpad�G?ٙ������labelspacing�G?�      �handlelength�G@       �handleheight�G?�ffffff�handletextpad�G?陙�����borderaxespad�G?�      �columnspacing�G@       �shadow��jvJ  K�_scatteryoffsets�hhK ��h��R�(KK��h!�C      �?�t�b�_legend_box�j�T  �VPacker���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�(j�T  j�T  �HPacker���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�j%U  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�(j3U  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�(j�T  �DrawingArea���)��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�j�T  ajU  h0h!C\����y@���R�h0h!C-؂-��{@���R����width�G@4      �height�G@      �xdescent�G        �ydescent�G        �_clip_children��jU  j�T  �dpi_transform�j�T  ubj�T  )��}�(j�7  j2T  h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�j2T  ajU  h0h!C@�~&f|@���R�h0h!C-؂-��{@���R���jU  j9T  jU  jBT  jU  �ubejU  h0h!C\����y@���R�h0h!C-؂-��{@���R���jnU  NjmU  N�sep�G@       �pad�K �mode��fixed��align�j�7  ubj3U  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�(jYU  )��}�(h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�j�T  ajU  h0h!C\����y@���R�h0h!C"""""Rz@���R���jmU  G@4      jnU  G@      joU  G        jpU  G        jqU  �jU  j�T  jrU  j�T  ubj�T  )��}�(j�7  j\T  h@�hANhBh>hChGhINhJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j2+  ]�j\T  ajU  h0h!C@�~&f|@���R�h0h!C"""""Rz@���R���jU  jaT  jU  jjT  jU  �ubejU  h0h!C\����y@���R�h0h!C"""""Rz@���R���jnU  NjmU  Nj�U  G@       j�U  K j�U  j�U  j�U  j�7  ubejU  h0h!C\����y@���R�h0h!C-؂-��{@���R���jnU  NjmU  Nj�U  G@      j�U  K j�U  j�U  j�U  j�7  ubajU  h0h!C\����y@���R�h0h!C-؂-��{@���R���jnU  NjmU  Nj�U  G@4      j�U  K j�U  j�U  j�U  j�7  ubejU  h�jT  �_findoffset���R�jnU  NjmU  Nj�U  G@      j�U  G@      j�U  j�U  j�U  j�7  ub�isaxes���parent�h>�_mode�N�_bbox_to_anchor�N�_shadow_props�}�(�ox�K�oy�J����u�legendPatch�j4+  �FancyBboxPatch���)��}�(h@�hANhBh>hChGhIjT  hJ�hK�hL�hMG?陙����hNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhl�hmNhnhohphs]�]�����hx�jI+  (G?陙����G?陙����G?陙����G?陙����t�jK+  �jL+  �0.8�jM+  j�U  jO+  jI  jV+  (G?�      G?�      G?�      G?陙����t�jX+  G?�333333jY+  K N��j[+  G        N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  j�  h0h!C���
�y@���R�j�  h0h!C�>�>�y@���R�js+  h0h!C���c@���R�jw+  h0h!C�`��K@���R��_bbox_transmuter�j4+  �BoxStyle.Round���)��}�(j�U  G        �rounding_size�G?ə�����ub�_mutation_scale�G@+�q�r�_mutation_aspect�Kub�
_alignment�j�7  �_legend_handle_box�j4U  �_loc_used_default���_outside_loc�N�	_loc_real�K �
_draggable�NubjYI  ]�j�I  �j�I  j�7  )��}�(h@�hANhBh>hChGhIjH  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  �$Residuals for LinearRegression Model�j�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�I  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  �center�j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�I  j�7  )��}�(h@�hANhBh>hChGhIjN  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G        j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�I  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j-7  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�I  j�7  )��}�(h@�hANhBh>hChGhIjQ  hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�j�  G?�      j�  G?�      j�7  hRj�6  j�7  j�7  j�7  )��}�(j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�I  j�7  j�7  j�7  Nj�7  G@(      j�7  j�7  ubj�7  �j�7  �j�7  �j�7  j�7  j�7  j�8  j�7  Nj�7  G        j�7  �j�7  Nj�7  Nj�7  G?�333333j�7  j�6  j_+  �ubj�I  jK  j�I  j6+  )��}�(h@�hANhBNhChGhIh�hJ�hK�hL�hMNhNNhONhP�hQhRhSNhT�hUNhV�hWhZ)��}�(h]]�h_ah`hbhc}�heK hfNhg��ubhiNhjNhkNhlNhmNhnhohphs]�]�����hx�jI+  jN+  jK+  �jL+  j7  jM+  jN+  jO+  jI  jV+  j�I  jX+  G        jY+  K N��j[+  K N��j]+  j^+  j_+  �j`+  Nja+  jg+  jh+  jm+  jn+  G        jo+  G        js+  G?�      jw+  G?�      j{+  G        j|+  j}+  j~+  G?�      ubj�I  �j�I  Nj�I  Nj�I  �j�I  Nj�I  }�h�]�(h�h>esj�I  Nubj+  Nj�7  Nj/I  Nj�I  N�colors�}�(�train_point�jK  �
test_point�j�T  j�E  j�6  u�hist���qqplot���_hax�h��_labels�]�(j�J  jKK  e�_colors�]�(jK  j�T  e�alphas�}�(jLV  G?�      jMV  G?�      u�train_score_�h0h!Cglk�T�?���R��test_score_�h0h!C�W�ע�?���R�ub.